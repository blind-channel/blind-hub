module raw_aes256(input w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, 
	output w50922, w50923, w50924, w50925, w50926, w50927, w50928, w50929, w50930, w50931, w50932, w50933, w50934, w50935, w50936, w50937, w50938, w50939, w50940, w50941, w50942, w50943, w50944, w50945, w50946, w50947, w50948, w50949, w50950, w50951, w50952, w50953, w50954, w50955, w50956, w50957, w50958, w50959, w50960, w50961, w50962, w50963, w50964, w50965, w50966, w50967, w50968, w50969, w50970, w50971, w50972, w50973, w50974, w50975, w50976, w50977, w50978, w50979, w50980, w50981, w50982, w50983, w50984, w50985, w50986, w50987, w50988, w50989, w50990, w50991, w50992, w50993, w50994, w50995, w50996, w50997, w50998, w50999, w51000, w51001, w51002, w51003, w51004, w51005, w51006, w51007, w51008, w51009, w51010, w51011, w51012, w51013, w51014, w51015, w51016, w51017, w51018, w51019, w51020, w51021, w51022, w51023, w51024, w51025, w51026, w51027, w51028, w51029, w51030, w51031, w51032, w51033, w51034, w51035, w51036, w51037, w51038, w51039, w51040, w51041, w51042, w51043, w51044, w51045, w51046, w51047, w51048, w51049);

	wire w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200, w19201, w19202, w19203, w19204, w19205, w19206, w19207, w19208, w19209, w19210, w19211, w19212, w19213, w19214, w19215, w19216, w19217, w19218, w19219, w19220, w19221, w19222, w19223, w19224, w19225, w19226, w19227, w19228, w19229, w19230, w19231, w19232, w19233, w19234, w19235, w19236, w19237, w19238, w19239, w19240, w19241, w19242, w19243, w19244, w19245, w19246, w19247, w19248, w19249, w19250, w19251, w19252, w19253, w19254, w19255, w19256, w19257, w19258, w19259, w19260, w19261, w19262, w19263, w19264, w19265, w19266, w19267, w19268, w19269, w19270, w19271, w19272, w19273, w19274, w19275, w19276, w19277, w19278, w19279, w19280, w19281, w19282, w19283, w19284, w19285, w19286, w19287, w19288, w19289, w19290, w19291, w19292, w19293, w19294, w19295, w19296, w19297, w19298, w19299, w19300, w19301, w19302, w19303, w19304, w19305, w19306, w19307, w19308, w19309, w19310, w19311, w19312, w19313, w19314, w19315, w19316, w19317, w19318, w19319, w19320, w19321, w19322, w19323, w19324, w19325, w19326, w19327, w19328, w19329, w19330, w19331, w19332, w19333, w19334, w19335, w19336, w19337, w19338, w19339, w19340, w19341, w19342, w19343, w19344, w19345, w19346, w19347, w19348, w19349, w19350, w19351, w19352, w19353, w19354, w19355, w19356, w19357, w19358, w19359, w19360, w19361, w19362, w19363, w19364, w19365, w19366, w19367, w19368, w19369, w19370, w19371, w19372, w19373, w19374, w19375, w19376, w19377, w19378, w19379, w19380, w19381, w19382, w19383, w19384, w19385, w19386, w19387, w19388, w19389, w19390, w19391, w19392, w19393, w19394, w19395, w19396, w19397, w19398, w19399, w19400, w19401, w19402, w19403, w19404, w19405, w19406, w19407, w19408, w19409, w19410, w19411, w19412, w19413, w19414, w19415, w19416, w19417, w19418, w19419, w19420, w19421, w19422, w19423, w19424, w19425, w19426, w19427, w19428, w19429, w19430, w19431, w19432, w19433, w19434, w19435, w19436, w19437, w19438, w19439, w19440, w19441, w19442, w19443, w19444, w19445, w19446, w19447, w19448, w19449, w19450, w19451, w19452, w19453, w19454, w19455, w19456, w19457, w19458, w19459, w19460, w19461, w19462, w19463, w19464, w19465, w19466, w19467, w19468, w19469, w19470, w19471, w19472, w19473, w19474, w19475, w19476, w19477, w19478, w19479, w19480, w19481, w19482, w19483, w19484, w19485, w19486, w19487, w19488, w19489, w19490, w19491, w19492, w19493, w19494, w19495, w19496, w19497, w19498, w19499, w19500, w19501, w19502, w19503, w19504, w19505, w19506, w19507, w19508, w19509, w19510, w19511, w19512, w19513, w19514, w19515, w19516, w19517, w19518, w19519, w19520, w19521, w19522, w19523, w19524, w19525, w19526, w19527, w19528, w19529, w19530, w19531, w19532, w19533, w19534, w19535, w19536, w19537, w19538, w19539, w19540, w19541, w19542, w19543, w19544, w19545, w19546, w19547, w19548, w19549, w19550, w19551, w19552, w19553, w19554, w19555, w19556, w19557, w19558, w19559, w19560, w19561, w19562, w19563, w19564, w19565, w19566, w19567, w19568, w19569, w19570, w19571, w19572, w19573, w19574, w19575, w19576, w19577, w19578, w19579, w19580, w19581, w19582, w19583, w19584, w19585, w19586, w19587, w19588, w19589, w19590, w19591, w19592, w19593, w19594, w19595, w19596, w19597, w19598, w19599, w19600, w19601, w19602, w19603, w19604, w19605, w19606, w19607, w19608, w19609, w19610, w19611, w19612, w19613, w19614, w19615, w19616, w19617, w19618, w19619, w19620, w19621, w19622, w19623, w19624, w19625, w19626, w19627, w19628, w19629, w19630, w19631, w19632, w19633, w19634, w19635, w19636, w19637, w19638, w19639, w19640, w19641, w19642, w19643, w19644, w19645, w19646, w19647, w19648, w19649, w19650, w19651, w19652, w19653, w19654, w19655, w19656, w19657, w19658, w19659, w19660, w19661, w19662, w19663, w19664, w19665, w19666, w19667, w19668, w19669, w19670, w19671, w19672, w19673, w19674, w19675, w19676, w19677, w19678, w19679, w19680, w19681, w19682, w19683, w19684, w19685, w19686, w19687, w19688, w19689, w19690, w19691, w19692, w19693, w19694, w19695, w19696, w19697, w19698, w19699, w19700, w19701, w19702, w19703, w19704, w19705, w19706, w19707, w19708, w19709, w19710, w19711, w19712, w19713, w19714, w19715, w19716, w19717, w19718, w19719, w19720, w19721, w19722, w19723, w19724, w19725, w19726, w19727, w19728, w19729, w19730, w19731, w19732, w19733, w19734, w19735, w19736, w19737, w19738, w19739, w19740, w19741, w19742, w19743, w19744, w19745, w19746, w19747, w19748, w19749, w19750, w19751, w19752, w19753, w19754, w19755, w19756, w19757, w19758, w19759, w19760, w19761, w19762, w19763, w19764, w19765, w19766, w19767, w19768, w19769, w19770, w19771, w19772, w19773, w19774, w19775, w19776, w19777, w19778, w19779, w19780, w19781, w19782, w19783, w19784, w19785, w19786, w19787, w19788, w19789, w19790, w19791, w19792, w19793, w19794, w19795, w19796, w19797, w19798, w19799, w19800, w19801, w19802, w19803, w19804, w19805, w19806, w19807, w19808, w19809, w19810, w19811, w19812, w19813, w19814, w19815, w19816, w19817, w19818, w19819, w19820, w19821, w19822, w19823, w19824, w19825, w19826, w19827, w19828, w19829, w19830, w19831, w19832, w19833, w19834, w19835, w19836, w19837, w19838, w19839, w19840, w19841, w19842, w19843, w19844, w19845, w19846, w19847, w19848, w19849, w19850, w19851, w19852, w19853, w19854, w19855, w19856, w19857, w19858, w19859, w19860, w19861, w19862, w19863, w19864, w19865, w19866, w19867, w19868, w19869, w19870, w19871, w19872, w19873, w19874, w19875, w19876, w19877, w19878, w19879, w19880, w19881, w19882, w19883, w19884, w19885, w19886, w19887, w19888, w19889, w19890, w19891, w19892, w19893, w19894, w19895, w19896, w19897, w19898, w19899, w19900, w19901, w19902, w19903, w19904, w19905, w19906, w19907, w19908, w19909, w19910, w19911, w19912, w19913, w19914, w19915, w19916, w19917, w19918, w19919, w19920, w19921, w19922, w19923, w19924, w19925, w19926, w19927, w19928, w19929, w19930, w19931, w19932, w19933, w19934, w19935, w19936, w19937, w19938, w19939, w19940, w19941, w19942, w19943, w19944, w19945, w19946, w19947, w19948, w19949, w19950, w19951, w19952, w19953, w19954, w19955, w19956, w19957, w19958, w19959, w19960, w19961, w19962, w19963, w19964, w19965, w19966, w19967, w19968, w19969, w19970, w19971, w19972, w19973, w19974, w19975, w19976, w19977, w19978, w19979, w19980, w19981, w19982, w19983, w19984, w19985, w19986, w19987, w19988, w19989, w19990, w19991, w19992, w19993, w19994, w19995, w19996, w19997, w19998, w19999, w20000, w20001, w20002, w20003, w20004, w20005, w20006, w20007, w20008, w20009, w20010, w20011, w20012, w20013, w20014, w20015, w20016, w20017, w20018, w20019, w20020, w20021, w20022, w20023, w20024, w20025, w20026, w20027, w20028, w20029, w20030, w20031, w20032, w20033, w20034, w20035, w20036, w20037, w20038, w20039, w20040, w20041, w20042, w20043, w20044, w20045, w20046, w20047, w20048, w20049, w20050, w20051, w20052, w20053, w20054, w20055, w20056, w20057, w20058, w20059, w20060, w20061, w20062, w20063, w20064, w20065, w20066, w20067, w20068, w20069, w20070, w20071, w20072, w20073, w20074, w20075, w20076, w20077, w20078, w20079, w20080, w20081, w20082, w20083, w20084, w20085, w20086, w20087, w20088, w20089, w20090, w20091, w20092, w20093, w20094, w20095, w20096, w20097, w20098, w20099, w20100, w20101, w20102, w20103, w20104, w20105, w20106, w20107, w20108, w20109, w20110, w20111, w20112, w20113, w20114, w20115, w20116, w20117, w20118, w20119, w20120, w20121, w20122, w20123, w20124, w20125, w20126, w20127, w20128, w20129, w20130, w20131, w20132, w20133, w20134, w20135, w20136, w20137, w20138, w20139, w20140, w20141, w20142, w20143, w20144, w20145, w20146, w20147, w20148, w20149, w20150, w20151, w20152, w20153, w20154, w20155, w20156, w20157, w20158, w20159, w20160, w20161, w20162, w20163, w20164, w20165, w20166, w20167, w20168, w20169, w20170, w20171, w20172, w20173, w20174, w20175, w20176, w20177, w20178, w20179, w20180, w20181, w20182, w20183, w20184, w20185, w20186, w20187, w20188, w20189, w20190, w20191, w20192, w20193, w20194, w20195, w20196, w20197, w20198, w20199, w20200, w20201, w20202, w20203, w20204, w20205, w20206, w20207, w20208, w20209, w20210, w20211, w20212, w20213, w20214, w20215, w20216, w20217, w20218, w20219, w20220, w20221, w20222, w20223, w20224, w20225, w20226, w20227, w20228, w20229, w20230, w20231, w20232, w20233, w20234, w20235, w20236, w20237, w20238, w20239, w20240, w20241, w20242, w20243, w20244, w20245, w20246, w20247, w20248, w20249, w20250, w20251, w20252, w20253, w20254, w20255, w20256, w20257, w20258, w20259, w20260, w20261, w20262, w20263, w20264, w20265, w20266, w20267, w20268, w20269, w20270, w20271, w20272, w20273, w20274, w20275, w20276, w20277, w20278, w20279, w20280, w20281, w20282, w20283, w20284, w20285, w20286, w20287, w20288, w20289, w20290, w20291, w20292, w20293, w20294, w20295, w20296, w20297, w20298, w20299, w20300, w20301, w20302, w20303, w20304, w20305, w20306, w20307, w20308, w20309, w20310, w20311, w20312, w20313, w20314, w20315, w20316, w20317, w20318, w20319, w20320, w20321, w20322, w20323, w20324, w20325, w20326, w20327, w20328, w20329, w20330, w20331, w20332, w20333, w20334, w20335, w20336, w20337, w20338, w20339, w20340, w20341, w20342, w20343, w20344, w20345, w20346, w20347, w20348, w20349, w20350, w20351, w20352, w20353, w20354, w20355, w20356, w20357, w20358, w20359, w20360, w20361, w20362, w20363, w20364, w20365, w20366, w20367, w20368, w20369, w20370, w20371, w20372, w20373, w20374, w20375, w20376, w20377, w20378, w20379, w20380, w20381, w20382, w20383, w20384, w20385, w20386, w20387, w20388, w20389, w20390, w20391, w20392, w20393, w20394, w20395, w20396, w20397, w20398, w20399, w20400, w20401, w20402, w20403, w20404, w20405, w20406, w20407, w20408, w20409, w20410, w20411, w20412, w20413, w20414, w20415, w20416, w20417, w20418, w20419, w20420, w20421, w20422, w20423, w20424, w20425, w20426, w20427, w20428, w20429, w20430, w20431, w20432, w20433, w20434, w20435, w20436, w20437, w20438, w20439, w20440, w20441, w20442, w20443, w20444, w20445, w20446, w20447, w20448, w20449, w20450, w20451, w20452, w20453, w20454, w20455, w20456, w20457, w20458, w20459, w20460, w20461, w20462, w20463, w20464, w20465, w20466, w20467, w20468, w20469, w20470, w20471, w20472, w20473, w20474, w20475, w20476, w20477, w20478, w20479, w20480, w20481, w20482, w20483, w20484, w20485, w20486, w20487, w20488, w20489, w20490, w20491, w20492, w20493, w20494, w20495, w20496, w20497, w20498, w20499, w20500, w20501, w20502, w20503, w20504, w20505, w20506, w20507, w20508, w20509, w20510, w20511, w20512, w20513, w20514, w20515, w20516, w20517, w20518, w20519, w20520, w20521, w20522, w20523, w20524, w20525, w20526, w20527, w20528, w20529, w20530, w20531, w20532, w20533, w20534, w20535, w20536, w20537, w20538, w20539, w20540, w20541, w20542, w20543, w20544, w20545, w20546, w20547, w20548, w20549, w20550, w20551, w20552, w20553, w20554, w20555, w20556, w20557, w20558, w20559, w20560, w20561, w20562, w20563, w20564, w20565, w20566, w20567, w20568, w20569, w20570, w20571, w20572, w20573, w20574, w20575, w20576, w20577, w20578, w20579, w20580, w20581, w20582, w20583, w20584, w20585, w20586, w20587, w20588, w20589, w20590, w20591, w20592, w20593, w20594, w20595, w20596, w20597, w20598, w20599, w20600, w20601, w20602, w20603, w20604, w20605, w20606, w20607, w20608, w20609, w20610, w20611, w20612, w20613, w20614, w20615, w20616, w20617, w20618, w20619, w20620, w20621, w20622, w20623, w20624, w20625, w20626, w20627, w20628, w20629, w20630, w20631, w20632, w20633, w20634, w20635, w20636, w20637, w20638, w20639, w20640, w20641, w20642, w20643, w20644, w20645, w20646, w20647, w20648, w20649, w20650, w20651, w20652, w20653, w20654, w20655, w20656, w20657, w20658, w20659, w20660, w20661, w20662, w20663, w20664, w20665, w20666, w20667, w20668, w20669, w20670, w20671, w20672, w20673, w20674, w20675, w20676, w20677, w20678, w20679, w20680, w20681, w20682, w20683, w20684, w20685, w20686, w20687, w20688, w20689, w20690, w20691, w20692, w20693, w20694, w20695, w20696, w20697, w20698, w20699, w20700, w20701, w20702, w20703, w20704, w20705, w20706, w20707, w20708, w20709, w20710, w20711, w20712, w20713, w20714, w20715, w20716, w20717, w20718, w20719, w20720, w20721, w20722, w20723, w20724, w20725, w20726, w20727, w20728, w20729, w20730, w20731, w20732, w20733, w20734, w20735, w20736, w20737, w20738, w20739, w20740, w20741, w20742, w20743, w20744, w20745, w20746, w20747, w20748, w20749, w20750, w20751, w20752, w20753, w20754, w20755, w20756, w20757, w20758, w20759, w20760, w20761, w20762, w20763, w20764, w20765, w20766, w20767, w20768, w20769, w20770, w20771, w20772, w20773, w20774, w20775, w20776, w20777, w20778, w20779, w20780, w20781, w20782, w20783, w20784, w20785, w20786, w20787, w20788, w20789, w20790, w20791, w20792, w20793, w20794, w20795, w20796, w20797, w20798, w20799, w20800, w20801, w20802, w20803, w20804, w20805, w20806, w20807, w20808, w20809, w20810, w20811, w20812, w20813, w20814, w20815, w20816, w20817, w20818, w20819, w20820, w20821, w20822, w20823, w20824, w20825, w20826, w20827, w20828, w20829, w20830, w20831, w20832, w20833, w20834, w20835, w20836, w20837, w20838, w20839, w20840, w20841, w20842, w20843, w20844, w20845, w20846, w20847, w20848, w20849, w20850, w20851, w20852, w20853, w20854, w20855, w20856, w20857, w20858, w20859, w20860, w20861, w20862, w20863, w20864, w20865, w20866, w20867, w20868, w20869, w20870, w20871, w20872, w20873, w20874, w20875, w20876, w20877, w20878, w20879, w20880, w20881, w20882, w20883, w20884, w20885, w20886, w20887, w20888, w20889, w20890, w20891, w20892, w20893, w20894, w20895, w20896, w20897, w20898, w20899, w20900, w20901, w20902, w20903, w20904, w20905, w20906, w20907, w20908, w20909, w20910, w20911, w20912, w20913, w20914, w20915, w20916, w20917, w20918, w20919, w20920, w20921, w20922, w20923, w20924, w20925, w20926, w20927, w20928, w20929, w20930, w20931, w20932, w20933, w20934, w20935, w20936, w20937, w20938, w20939, w20940, w20941, w20942, w20943, w20944, w20945, w20946, w20947, w20948, w20949, w20950, w20951, w20952, w20953, w20954, w20955, w20956, w20957, w20958, w20959, w20960, w20961, w20962, w20963, w20964, w20965, w20966, w20967, w20968, w20969, w20970, w20971, w20972, w20973, w20974, w20975, w20976, w20977, w20978, w20979, w20980, w20981, w20982, w20983, w20984, w20985, w20986, w20987, w20988, w20989, w20990, w20991, w20992, w20993, w20994, w20995, w20996, w20997, w20998, w20999, w21000, w21001, w21002, w21003, w21004, w21005, w21006, w21007, w21008, w21009, w21010, w21011, w21012, w21013, w21014, w21015, w21016, w21017, w21018, w21019, w21020, w21021, w21022, w21023, w21024, w21025, w21026, w21027, w21028, w21029, w21030, w21031, w21032, w21033, w21034, w21035, w21036, w21037, w21038, w21039, w21040, w21041, w21042, w21043, w21044, w21045, w21046, w21047, w21048, w21049, w21050, w21051, w21052, w21053, w21054, w21055, w21056, w21057, w21058, w21059, w21060, w21061, w21062, w21063, w21064, w21065, w21066, w21067, w21068, w21069, w21070, w21071, w21072, w21073, w21074, w21075, w21076, w21077, w21078, w21079, w21080, w21081, w21082, w21083, w21084, w21085, w21086, w21087, w21088, w21089, w21090, w21091, w21092, w21093, w21094, w21095, w21096, w21097, w21098, w21099, w21100, w21101, w21102, w21103, w21104, w21105, w21106, w21107, w21108, w21109, w21110, w21111, w21112, w21113, w21114, w21115, w21116, w21117, w21118, w21119, w21120, w21121, w21122, w21123, w21124, w21125, w21126, w21127, w21128, w21129, w21130, w21131, w21132, w21133, w21134, w21135, w21136, w21137, w21138, w21139, w21140, w21141, w21142, w21143, w21144, w21145, w21146, w21147, w21148, w21149, w21150, w21151, w21152, w21153, w21154, w21155, w21156, w21157, w21158, w21159, w21160, w21161, w21162, w21163, w21164, w21165, w21166, w21167, w21168, w21169, w21170, w21171, w21172, w21173, w21174, w21175, w21176, w21177, w21178, w21179, w21180, w21181, w21182, w21183, w21184, w21185, w21186, w21187, w21188, w21189, w21190, w21191, w21192, w21193, w21194, w21195, w21196, w21197, w21198, w21199, w21200, w21201, w21202, w21203, w21204, w21205, w21206, w21207, w21208, w21209, w21210, w21211, w21212, w21213, w21214, w21215, w21216, w21217, w21218, w21219, w21220, w21221, w21222, w21223, w21224, w21225, w21226, w21227, w21228, w21229, w21230, w21231, w21232, w21233, w21234, w21235, w21236, w21237, w21238, w21239, w21240, w21241, w21242, w21243, w21244, w21245, w21246, w21247, w21248, w21249, w21250, w21251, w21252, w21253, w21254, w21255, w21256, w21257, w21258, w21259, w21260, w21261, w21262, w21263, w21264, w21265, w21266, w21267, w21268, w21269, w21270, w21271, w21272, w21273, w21274, w21275, w21276, w21277, w21278, w21279, w21280, w21281, w21282, w21283, w21284, w21285, w21286, w21287, w21288, w21289, w21290, w21291, w21292, w21293, w21294, w21295, w21296, w21297, w21298, w21299, w21300, w21301, w21302, w21303, w21304, w21305, w21306, w21307, w21308, w21309, w21310, w21311, w21312, w21313, w21314, w21315, w21316, w21317, w21318, w21319, w21320, w21321, w21322, w21323, w21324, w21325, w21326, w21327, w21328, w21329, w21330, w21331, w21332, w21333, w21334, w21335, w21336, w21337, w21338, w21339, w21340, w21341, w21342, w21343, w21344, w21345, w21346, w21347, w21348, w21349, w21350, w21351, w21352, w21353, w21354, w21355, w21356, w21357, w21358, w21359, w21360, w21361, w21362, w21363, w21364, w21365, w21366, w21367, w21368, w21369, w21370, w21371, w21372, w21373, w21374, w21375, w21376, w21377, w21378, w21379, w21380, w21381, w21382, w21383, w21384, w21385, w21386, w21387, w21388, w21389, w21390, w21391, w21392, w21393, w21394, w21395, w21396, w21397, w21398, w21399, w21400, w21401, w21402, w21403, w21404, w21405, w21406, w21407, w21408, w21409, w21410, w21411, w21412, w21413, w21414, w21415, w21416, w21417, w21418, w21419, w21420, w21421, w21422, w21423, w21424, w21425, w21426, w21427, w21428, w21429, w21430, w21431, w21432, w21433, w21434, w21435, w21436, w21437, w21438, w21439, w21440, w21441, w21442, w21443, w21444, w21445, w21446, w21447, w21448, w21449, w21450, w21451, w21452, w21453, w21454, w21455, w21456, w21457, w21458, w21459, w21460, w21461, w21462, w21463, w21464, w21465, w21466, w21467, w21468, w21469, w21470, w21471, w21472, w21473, w21474, w21475, w21476, w21477, w21478, w21479, w21480, w21481, w21482, w21483, w21484, w21485, w21486, w21487, w21488, w21489, w21490, w21491, w21492, w21493, w21494, w21495, w21496, w21497, w21498, w21499, w21500, w21501, w21502, w21503, w21504, w21505, w21506, w21507, w21508, w21509, w21510, w21511, w21512, w21513, w21514, w21515, w21516, w21517, w21518, w21519, w21520, w21521, w21522, w21523, w21524, w21525, w21526, w21527, w21528, w21529, w21530, w21531, w21532, w21533, w21534, w21535, w21536, w21537, w21538, w21539, w21540, w21541, w21542, w21543, w21544, w21545, w21546, w21547, w21548, w21549, w21550, w21551, w21552, w21553, w21554, w21555, w21556, w21557, w21558, w21559, w21560, w21561, w21562, w21563, w21564, w21565, w21566, w21567, w21568, w21569, w21570, w21571, w21572, w21573, w21574, w21575, w21576, w21577, w21578, w21579, w21580, w21581, w21582, w21583, w21584, w21585, w21586, w21587, w21588, w21589, w21590, w21591, w21592, w21593, w21594, w21595, w21596, w21597, w21598, w21599, w21600, w21601, w21602, w21603, w21604, w21605, w21606, w21607, w21608, w21609, w21610, w21611, w21612, w21613, w21614, w21615, w21616, w21617, w21618, w21619, w21620, w21621, w21622, w21623, w21624, w21625, w21626, w21627, w21628, w21629, w21630, w21631, w21632, w21633, w21634, w21635, w21636, w21637, w21638, w21639, w21640, w21641, w21642, w21643, w21644, w21645, w21646, w21647, w21648, w21649, w21650, w21651, w21652, w21653, w21654, w21655, w21656, w21657, w21658, w21659, w21660, w21661, w21662, w21663, w21664, w21665, w21666, w21667, w21668, w21669, w21670, w21671, w21672, w21673, w21674, w21675, w21676, w21677, w21678, w21679, w21680, w21681, w21682, w21683, w21684, w21685, w21686, w21687, w21688, w21689, w21690, w21691, w21692, w21693, w21694, w21695, w21696, w21697, w21698, w21699, w21700, w21701, w21702, w21703, w21704, w21705, w21706, w21707, w21708, w21709, w21710, w21711, w21712, w21713, w21714, w21715, w21716, w21717, w21718, w21719, w21720, w21721, w21722, w21723, w21724, w21725, w21726, w21727, w21728, w21729, w21730, w21731, w21732, w21733, w21734, w21735, w21736, w21737, w21738, w21739, w21740, w21741, w21742, w21743, w21744, w21745, w21746, w21747, w21748, w21749, w21750, w21751, w21752, w21753, w21754, w21755, w21756, w21757, w21758, w21759, w21760, w21761, w21762, w21763, w21764, w21765, w21766, w21767, w21768, w21769, w21770, w21771, w21772, w21773, w21774, w21775, w21776, w21777, w21778, w21779, w21780, w21781, w21782, w21783, w21784, w21785, w21786, w21787, w21788, w21789, w21790, w21791, w21792, w21793, w21794, w21795, w21796, w21797, w21798, w21799, w21800, w21801, w21802, w21803, w21804, w21805, w21806, w21807, w21808, w21809, w21810, w21811, w21812, w21813, w21814, w21815, w21816, w21817, w21818, w21819, w21820, w21821, w21822, w21823, w21824, w21825, w21826, w21827, w21828, w21829, w21830, w21831, w21832, w21833, w21834, w21835, w21836, w21837, w21838, w21839, w21840, w21841, w21842, w21843, w21844, w21845, w21846, w21847, w21848, w21849, w21850, w21851, w21852, w21853, w21854, w21855, w21856, w21857, w21858, w21859, w21860, w21861, w21862, w21863, w21864, w21865, w21866, w21867, w21868, w21869, w21870, w21871, w21872, w21873, w21874, w21875, w21876, w21877, w21878, w21879, w21880, w21881, w21882, w21883, w21884, w21885, w21886, w21887, w21888, w21889, w21890, w21891, w21892, w21893, w21894, w21895, w21896, w21897, w21898, w21899, w21900, w21901, w21902, w21903, w21904, w21905, w21906, w21907, w21908, w21909, w21910, w21911, w21912, w21913, w21914, w21915, w21916, w21917, w21918, w21919, w21920, w21921, w21922, w21923, w21924, w21925, w21926, w21927, w21928, w21929, w21930, w21931, w21932, w21933, w21934, w21935, w21936, w21937, w21938, w21939, w21940, w21941, w21942, w21943, w21944, w21945, w21946, w21947, w21948, w21949, w21950, w21951, w21952, w21953, w21954, w21955, w21956, w21957, w21958, w21959, w21960, w21961, w21962, w21963, w21964, w21965, w21966, w21967, w21968, w21969, w21970, w21971, w21972, w21973, w21974, w21975, w21976, w21977, w21978, w21979, w21980, w21981, w21982, w21983, w21984, w21985, w21986, w21987, w21988, w21989, w21990, w21991, w21992, w21993, w21994, w21995, w21996, w21997, w21998, w21999, w22000, w22001, w22002, w22003, w22004, w22005, w22006, w22007, w22008, w22009, w22010, w22011, w22012, w22013, w22014, w22015, w22016, w22017, w22018, w22019, w22020, w22021, w22022, w22023, w22024, w22025, w22026, w22027, w22028, w22029, w22030, w22031, w22032, w22033, w22034, w22035, w22036, w22037, w22038, w22039, w22040, w22041, w22042, w22043, w22044, w22045, w22046, w22047, w22048, w22049, w22050, w22051, w22052, w22053, w22054, w22055, w22056, w22057, w22058, w22059, w22060, w22061, w22062, w22063, w22064, w22065, w22066, w22067, w22068, w22069, w22070, w22071, w22072, w22073, w22074, w22075, w22076, w22077, w22078, w22079, w22080, w22081, w22082, w22083, w22084, w22085, w22086, w22087, w22088, w22089, w22090, w22091, w22092, w22093, w22094, w22095, w22096, w22097, w22098, w22099, w22100, w22101, w22102, w22103, w22104, w22105, w22106, w22107, w22108, w22109, w22110, w22111, w22112, w22113, w22114, w22115, w22116, w22117, w22118, w22119, w22120, w22121, w22122, w22123, w22124, w22125, w22126, w22127, w22128, w22129, w22130, w22131, w22132, w22133, w22134, w22135, w22136, w22137, w22138, w22139, w22140, w22141, w22142, w22143, w22144, w22145, w22146, w22147, w22148, w22149, w22150, w22151, w22152, w22153, w22154, w22155, w22156, w22157, w22158, w22159, w22160, w22161, w22162, w22163, w22164, w22165, w22166, w22167, w22168, w22169, w22170, w22171, w22172, w22173, w22174, w22175, w22176, w22177, w22178, w22179, w22180, w22181, w22182, w22183, w22184, w22185, w22186, w22187, w22188, w22189, w22190, w22191, w22192, w22193, w22194, w22195, w22196, w22197, w22198, w22199, w22200, w22201, w22202, w22203, w22204, w22205, w22206, w22207, w22208, w22209, w22210, w22211, w22212, w22213, w22214, w22215, w22216, w22217, w22218, w22219, w22220, w22221, w22222, w22223, w22224, w22225, w22226, w22227, w22228, w22229, w22230, w22231, w22232, w22233, w22234, w22235, w22236, w22237, w22238, w22239, w22240, w22241, w22242, w22243, w22244, w22245, w22246, w22247, w22248, w22249, w22250, w22251, w22252, w22253, w22254, w22255, w22256, w22257, w22258, w22259, w22260, w22261, w22262, w22263, w22264, w22265, w22266, w22267, w22268, w22269, w22270, w22271, w22272, w22273, w22274, w22275, w22276, w22277, w22278, w22279, w22280, w22281, w22282, w22283, w22284, w22285, w22286, w22287, w22288, w22289, w22290, w22291, w22292, w22293, w22294, w22295, w22296, w22297, w22298, w22299, w22300, w22301, w22302, w22303, w22304, w22305, w22306, w22307, w22308, w22309, w22310, w22311, w22312, w22313, w22314, w22315, w22316, w22317, w22318, w22319, w22320, w22321, w22322, w22323, w22324, w22325, w22326, w22327, w22328, w22329, w22330, w22331, w22332, w22333, w22334, w22335, w22336, w22337, w22338, w22339, w22340, w22341, w22342, w22343, w22344, w22345, w22346, w22347, w22348, w22349, w22350, w22351, w22352, w22353, w22354, w22355, w22356, w22357, w22358, w22359, w22360, w22361, w22362, w22363, w22364, w22365, w22366, w22367, w22368, w22369, w22370, w22371, w22372, w22373, w22374, w22375, w22376, w22377, w22378, w22379, w22380, w22381, w22382, w22383, w22384, w22385, w22386, w22387, w22388, w22389, w22390, w22391, w22392, w22393, w22394, w22395, w22396, w22397, w22398, w22399, w22400, w22401, w22402, w22403, w22404, w22405, w22406, w22407, w22408, w22409, w22410, w22411, w22412, w22413, w22414, w22415, w22416, w22417, w22418, w22419, w22420, w22421, w22422, w22423, w22424, w22425, w22426, w22427, w22428, w22429, w22430, w22431, w22432, w22433, w22434, w22435, w22436, w22437, w22438, w22439, w22440, w22441, w22442, w22443, w22444, w22445, w22446, w22447, w22448, w22449, w22450, w22451, w22452, w22453, w22454, w22455, w22456, w22457, w22458, w22459, w22460, w22461, w22462, w22463, w22464, w22465, w22466, w22467, w22468, w22469, w22470, w22471, w22472, w22473, w22474, w22475, w22476, w22477, w22478, w22479, w22480, w22481, w22482, w22483, w22484, w22485, w22486, w22487, w22488, w22489, w22490, w22491, w22492, w22493, w22494, w22495, w22496, w22497, w22498, w22499, w22500, w22501, w22502, w22503, w22504, w22505, w22506, w22507, w22508, w22509, w22510, w22511, w22512, w22513, w22514, w22515, w22516, w22517, w22518, w22519, w22520, w22521, w22522, w22523, w22524, w22525, w22526, w22527, w22528, w22529, w22530, w22531, w22532, w22533, w22534, w22535, w22536, w22537, w22538, w22539, w22540, w22541, w22542, w22543, w22544, w22545, w22546, w22547, w22548, w22549, w22550, w22551, w22552, w22553, w22554, w22555, w22556, w22557, w22558, w22559, w22560, w22561, w22562, w22563, w22564, w22565, w22566, w22567, w22568, w22569, w22570, w22571, w22572, w22573, w22574, w22575, w22576, w22577, w22578, w22579, w22580, w22581, w22582, w22583, w22584, w22585, w22586, w22587, w22588, w22589, w22590, w22591, w22592, w22593, w22594, w22595, w22596, w22597, w22598, w22599, w22600, w22601, w22602, w22603, w22604, w22605, w22606, w22607, w22608, w22609, w22610, w22611, w22612, w22613, w22614, w22615, w22616, w22617, w22618, w22619, w22620, w22621, w22622, w22623, w22624, w22625, w22626, w22627, w22628, w22629, w22630, w22631, w22632, w22633, w22634, w22635, w22636, w22637, w22638, w22639, w22640, w22641, w22642, w22643, w22644, w22645, w22646, w22647, w22648, w22649, w22650, w22651, w22652, w22653, w22654, w22655, w22656, w22657, w22658, w22659, w22660, w22661, w22662, w22663, w22664, w22665, w22666, w22667, w22668, w22669, w22670, w22671, w22672, w22673, w22674, w22675, w22676, w22677, w22678, w22679, w22680, w22681, w22682, w22683, w22684, w22685, w22686, w22687, w22688, w22689, w22690, w22691, w22692, w22693, w22694, w22695, w22696, w22697, w22698, w22699, w22700, w22701, w22702, w22703, w22704, w22705, w22706, w22707, w22708, w22709, w22710, w22711, w22712, w22713, w22714, w22715, w22716, w22717, w22718, w22719, w22720, w22721, w22722, w22723, w22724, w22725, w22726, w22727, w22728, w22729, w22730, w22731, w22732, w22733, w22734, w22735, w22736, w22737, w22738, w22739, w22740, w22741, w22742, w22743, w22744, w22745, w22746, w22747, w22748, w22749, w22750, w22751, w22752, w22753, w22754, w22755, w22756, w22757, w22758, w22759, w22760, w22761, w22762, w22763, w22764, w22765, w22766, w22767, w22768, w22769, w22770, w22771, w22772, w22773, w22774, w22775, w22776, w22777, w22778, w22779, w22780, w22781, w22782, w22783, w22784, w22785, w22786, w22787, w22788, w22789, w22790, w22791, w22792, w22793, w22794, w22795, w22796, w22797, w22798, w22799, w22800, w22801, w22802, w22803, w22804, w22805, w22806, w22807, w22808, w22809, w22810, w22811, w22812, w22813, w22814, w22815, w22816, w22817, w22818, w22819, w22820, w22821, w22822, w22823, w22824, w22825, w22826, w22827, w22828, w22829, w22830, w22831, w22832, w22833, w22834, w22835, w22836, w22837, w22838, w22839, w22840, w22841, w22842, w22843, w22844, w22845, w22846, w22847, w22848, w22849, w22850, w22851, w22852, w22853, w22854, w22855, w22856, w22857, w22858, w22859, w22860, w22861, w22862, w22863, w22864, w22865, w22866, w22867, w22868, w22869, w22870, w22871, w22872, w22873, w22874, w22875, w22876, w22877, w22878, w22879, w22880, w22881, w22882, w22883, w22884, w22885, w22886, w22887, w22888, w22889, w22890, w22891, w22892, w22893, w22894, w22895, w22896, w22897, w22898, w22899, w22900, w22901, w22902, w22903, w22904, w22905, w22906, w22907, w22908, w22909, w22910, w22911, w22912, w22913, w22914, w22915, w22916, w22917, w22918, w22919, w22920, w22921, w22922, w22923, w22924, w22925, w22926, w22927, w22928, w22929, w22930, w22931, w22932, w22933, w22934, w22935, w22936, w22937, w22938, w22939, w22940, w22941, w22942, w22943, w22944, w22945, w22946, w22947, w22948, w22949, w22950, w22951, w22952, w22953, w22954, w22955, w22956, w22957, w22958, w22959, w22960, w22961, w22962, w22963, w22964, w22965, w22966, w22967, w22968, w22969, w22970, w22971, w22972, w22973, w22974, w22975, w22976, w22977, w22978, w22979, w22980, w22981, w22982, w22983, w22984, w22985, w22986, w22987, w22988, w22989, w22990, w22991, w22992, w22993, w22994, w22995, w22996, w22997, w22998, w22999, w23000, w23001, w23002, w23003, w23004, w23005, w23006, w23007, w23008, w23009, w23010, w23011, w23012, w23013, w23014, w23015, w23016, w23017, w23018, w23019, w23020, w23021, w23022, w23023, w23024, w23025, w23026, w23027, w23028, w23029, w23030, w23031, w23032, w23033, w23034, w23035, w23036, w23037, w23038, w23039, w23040, w23041, w23042, w23043, w23044, w23045, w23046, w23047, w23048, w23049, w23050, w23051, w23052, w23053, w23054, w23055, w23056, w23057, w23058, w23059, w23060, w23061, w23062, w23063, w23064, w23065, w23066, w23067, w23068, w23069, w23070, w23071, w23072, w23073, w23074, w23075, w23076, w23077, w23078, w23079, w23080, w23081, w23082, w23083, w23084, w23085, w23086, w23087, w23088, w23089, w23090, w23091, w23092, w23093, w23094, w23095, w23096, w23097, w23098, w23099, w23100, w23101, w23102, w23103, w23104, w23105, w23106, w23107, w23108, w23109, w23110, w23111, w23112, w23113, w23114, w23115, w23116, w23117, w23118, w23119, w23120, w23121, w23122, w23123, w23124, w23125, w23126, w23127, w23128, w23129, w23130, w23131, w23132, w23133, w23134, w23135, w23136, w23137, w23138, w23139, w23140, w23141, w23142, w23143, w23144, w23145, w23146, w23147, w23148, w23149, w23150, w23151, w23152, w23153, w23154, w23155, w23156, w23157, w23158, w23159, w23160, w23161, w23162, w23163, w23164, w23165, w23166, w23167, w23168, w23169, w23170, w23171, w23172, w23173, w23174, w23175, w23176, w23177, w23178, w23179, w23180, w23181, w23182, w23183, w23184, w23185, w23186, w23187, w23188, w23189, w23190, w23191, w23192, w23193, w23194, w23195, w23196, w23197, w23198, w23199, w23200, w23201, w23202, w23203, w23204, w23205, w23206, w23207, w23208, w23209, w23210, w23211, w23212, w23213, w23214, w23215, w23216, w23217, w23218, w23219, w23220, w23221, w23222, w23223, w23224, w23225, w23226, w23227, w23228, w23229, w23230, w23231, w23232, w23233, w23234, w23235, w23236, w23237, w23238, w23239, w23240, w23241, w23242, w23243, w23244, w23245, w23246, w23247, w23248, w23249, w23250, w23251, w23252, w23253, w23254, w23255, w23256, w23257, w23258, w23259, w23260, w23261, w23262, w23263, w23264, w23265, w23266, w23267, w23268, w23269, w23270, w23271, w23272, w23273, w23274, w23275, w23276, w23277, w23278, w23279, w23280, w23281, w23282, w23283, w23284, w23285, w23286, w23287, w23288, w23289, w23290, w23291, w23292, w23293, w23294, w23295, w23296, w23297, w23298, w23299, w23300, w23301, w23302, w23303, w23304, w23305, w23306, w23307, w23308, w23309, w23310, w23311, w23312, w23313, w23314, w23315, w23316, w23317, w23318, w23319, w23320, w23321, w23322, w23323, w23324, w23325, w23326, w23327, w23328, w23329, w23330, w23331, w23332, w23333, w23334, w23335, w23336, w23337, w23338, w23339, w23340, w23341, w23342, w23343, w23344, w23345, w23346, w23347, w23348, w23349, w23350, w23351, w23352, w23353, w23354, w23355, w23356, w23357, w23358, w23359, w23360, w23361, w23362, w23363, w23364, w23365, w23366, w23367, w23368, w23369, w23370, w23371, w23372, w23373, w23374, w23375, w23376, w23377, w23378, w23379, w23380, w23381, w23382, w23383, w23384, w23385, w23386, w23387, w23388, w23389, w23390, w23391, w23392, w23393, w23394, w23395, w23396, w23397, w23398, w23399, w23400, w23401, w23402, w23403, w23404, w23405, w23406, w23407, w23408, w23409, w23410, w23411, w23412, w23413, w23414, w23415, w23416, w23417, w23418, w23419, w23420, w23421, w23422, w23423, w23424, w23425, w23426, w23427, w23428, w23429, w23430, w23431, w23432, w23433, w23434, w23435, w23436, w23437, w23438, w23439, w23440, w23441, w23442, w23443, w23444, w23445, w23446, w23447, w23448, w23449, w23450, w23451, w23452, w23453, w23454, w23455, w23456, w23457, w23458, w23459, w23460, w23461, w23462, w23463, w23464, w23465, w23466, w23467, w23468, w23469, w23470, w23471, w23472, w23473, w23474, w23475, w23476, w23477, w23478, w23479, w23480, w23481, w23482, w23483, w23484, w23485, w23486, w23487, w23488, w23489, w23490, w23491, w23492, w23493, w23494, w23495, w23496, w23497, w23498, w23499, w23500, w23501, w23502, w23503, w23504, w23505, w23506, w23507, w23508, w23509, w23510, w23511, w23512, w23513, w23514, w23515, w23516, w23517, w23518, w23519, w23520, w23521, w23522, w23523, w23524, w23525, w23526, w23527, w23528, w23529, w23530, w23531, w23532, w23533, w23534, w23535, w23536, w23537, w23538, w23539, w23540, w23541, w23542, w23543, w23544, w23545, w23546, w23547, w23548, w23549, w23550, w23551, w23552, w23553, w23554, w23555, w23556, w23557, w23558, w23559, w23560, w23561, w23562, w23563, w23564, w23565, w23566, w23567, w23568, w23569, w23570, w23571, w23572, w23573, w23574, w23575, w23576, w23577, w23578, w23579, w23580, w23581, w23582, w23583, w23584, w23585, w23586, w23587, w23588, w23589, w23590, w23591, w23592, w23593, w23594, w23595, w23596, w23597, w23598, w23599, w23600, w23601, w23602, w23603, w23604, w23605, w23606, w23607, w23608, w23609, w23610, w23611, w23612, w23613, w23614, w23615, w23616, w23617, w23618, w23619, w23620, w23621, w23622, w23623, w23624, w23625, w23626, w23627, w23628, w23629, w23630, w23631, w23632, w23633, w23634, w23635, w23636, w23637, w23638, w23639, w23640, w23641, w23642, w23643, w23644, w23645, w23646, w23647, w23648, w23649, w23650, w23651, w23652, w23653, w23654, w23655, w23656, w23657, w23658, w23659, w23660, w23661, w23662, w23663, w23664, w23665, w23666, w23667, w23668, w23669, w23670, w23671, w23672, w23673, w23674, w23675, w23676, w23677, w23678, w23679, w23680, w23681, w23682, w23683, w23684, w23685, w23686, w23687, w23688, w23689, w23690, w23691, w23692, w23693, w23694, w23695, w23696, w23697, w23698, w23699, w23700, w23701, w23702, w23703, w23704, w23705, w23706, w23707, w23708, w23709, w23710, w23711, w23712, w23713, w23714, w23715, w23716, w23717, w23718, w23719, w23720, w23721, w23722, w23723, w23724, w23725, w23726, w23727, w23728, w23729, w23730, w23731, w23732, w23733, w23734, w23735, w23736, w23737, w23738, w23739, w23740, w23741, w23742, w23743, w23744, w23745, w23746, w23747, w23748, w23749, w23750, w23751, w23752, w23753, w23754, w23755, w23756, w23757, w23758, w23759, w23760, w23761, w23762, w23763, w23764, w23765, w23766, w23767, w23768, w23769, w23770, w23771, w23772, w23773, w23774, w23775, w23776, w23777, w23778, w23779, w23780, w23781, w23782, w23783, w23784, w23785, w23786, w23787, w23788, w23789, w23790, w23791, w23792, w23793, w23794, w23795, w23796, w23797, w23798, w23799, w23800, w23801, w23802, w23803, w23804, w23805, w23806, w23807, w23808, w23809, w23810, w23811, w23812, w23813, w23814, w23815, w23816, w23817, w23818, w23819, w23820, w23821, w23822, w23823, w23824, w23825, w23826, w23827, w23828, w23829, w23830, w23831, w23832, w23833, w23834, w23835, w23836, w23837, w23838, w23839, w23840, w23841, w23842, w23843, w23844, w23845, w23846, w23847, w23848, w23849, w23850, w23851, w23852, w23853, w23854, w23855, w23856, w23857, w23858, w23859, w23860, w23861, w23862, w23863, w23864, w23865, w23866, w23867, w23868, w23869, w23870, w23871, w23872, w23873, w23874, w23875, w23876, w23877, w23878, w23879, w23880, w23881, w23882, w23883, w23884, w23885, w23886, w23887, w23888, w23889, w23890, w23891, w23892, w23893, w23894, w23895, w23896, w23897, w23898, w23899, w23900, w23901, w23902, w23903, w23904, w23905, w23906, w23907, w23908, w23909, w23910, w23911, w23912, w23913, w23914, w23915, w23916, w23917, w23918, w23919, w23920, w23921, w23922, w23923, w23924, w23925, w23926, w23927, w23928, w23929, w23930, w23931, w23932, w23933, w23934, w23935, w23936, w23937, w23938, w23939, w23940, w23941, w23942, w23943, w23944, w23945, w23946, w23947, w23948, w23949, w23950, w23951, w23952, w23953, w23954, w23955, w23956, w23957, w23958, w23959, w23960, w23961, w23962, w23963, w23964, w23965, w23966, w23967, w23968, w23969, w23970, w23971, w23972, w23973, w23974, w23975, w23976, w23977, w23978, w23979, w23980, w23981, w23982, w23983, w23984, w23985, w23986, w23987, w23988, w23989, w23990, w23991, w23992, w23993, w23994, w23995, w23996, w23997, w23998, w23999, w24000, w24001, w24002, w24003, w24004, w24005, w24006, w24007, w24008, w24009, w24010, w24011, w24012, w24013, w24014, w24015, w24016, w24017, w24018, w24019, w24020, w24021, w24022, w24023, w24024, w24025, w24026, w24027, w24028, w24029, w24030, w24031, w24032, w24033, w24034, w24035, w24036, w24037, w24038, w24039, w24040, w24041, w24042, w24043, w24044, w24045, w24046, w24047, w24048, w24049, w24050, w24051, w24052, w24053, w24054, w24055, w24056, w24057, w24058, w24059, w24060, w24061, w24062, w24063, w24064, w24065, w24066, w24067, w24068, w24069, w24070, w24071, w24072, w24073, w24074, w24075, w24076, w24077, w24078, w24079, w24080, w24081, w24082, w24083, w24084, w24085, w24086, w24087, w24088, w24089, w24090, w24091, w24092, w24093, w24094, w24095, w24096, w24097, w24098, w24099, w24100, w24101, w24102, w24103, w24104, w24105, w24106, w24107, w24108, w24109, w24110, w24111, w24112, w24113, w24114, w24115, w24116, w24117, w24118, w24119, w24120, w24121, w24122, w24123, w24124, w24125, w24126, w24127, w24128, w24129, w24130, w24131, w24132, w24133, w24134, w24135, w24136, w24137, w24138, w24139, w24140, w24141, w24142, w24143, w24144, w24145, w24146, w24147, w24148, w24149, w24150, w24151, w24152, w24153, w24154, w24155, w24156, w24157, w24158, w24159, w24160, w24161, w24162, w24163, w24164, w24165, w24166, w24167, w24168, w24169, w24170, w24171, w24172, w24173, w24174, w24175, w24176, w24177, w24178, w24179, w24180, w24181, w24182, w24183, w24184, w24185, w24186, w24187, w24188, w24189, w24190, w24191, w24192, w24193, w24194, w24195, w24196, w24197, w24198, w24199, w24200, w24201, w24202, w24203, w24204, w24205, w24206, w24207, w24208, w24209, w24210, w24211, w24212, w24213, w24214, w24215, w24216, w24217, w24218, w24219, w24220, w24221, w24222, w24223, w24224, w24225, w24226, w24227, w24228, w24229, w24230, w24231, w24232, w24233, w24234, w24235, w24236, w24237, w24238, w24239, w24240, w24241, w24242, w24243, w24244, w24245, w24246, w24247, w24248, w24249, w24250, w24251, w24252, w24253, w24254, w24255, w24256, w24257, w24258, w24259, w24260, w24261, w24262, w24263, w24264, w24265, w24266, w24267, w24268, w24269, w24270, w24271, w24272, w24273, w24274, w24275, w24276, w24277, w24278, w24279, w24280, w24281, w24282, w24283, w24284, w24285, w24286, w24287, w24288, w24289, w24290, w24291, w24292, w24293, w24294, w24295, w24296, w24297, w24298, w24299, w24300, w24301, w24302, w24303, w24304, w24305, w24306, w24307, w24308, w24309, w24310, w24311, w24312, w24313, w24314, w24315, w24316, w24317, w24318, w24319, w24320, w24321, w24322, w24323, w24324, w24325, w24326, w24327, w24328, w24329, w24330, w24331, w24332, w24333, w24334, w24335, w24336, w24337, w24338, w24339, w24340, w24341, w24342, w24343, w24344, w24345, w24346, w24347, w24348, w24349, w24350, w24351, w24352, w24353, w24354, w24355, w24356, w24357, w24358, w24359, w24360, w24361, w24362, w24363, w24364, w24365, w24366, w24367, w24368, w24369, w24370, w24371, w24372, w24373, w24374, w24375, w24376, w24377, w24378, w24379, w24380, w24381, w24382, w24383, w24384, w24385, w24386, w24387, w24388, w24389, w24390, w24391, w24392, w24393, w24394, w24395, w24396, w24397, w24398, w24399, w24400, w24401, w24402, w24403, w24404, w24405, w24406, w24407, w24408, w24409, w24410, w24411, w24412, w24413, w24414, w24415, w24416, w24417, w24418, w24419, w24420, w24421, w24422, w24423, w24424, w24425, w24426, w24427, w24428, w24429, w24430, w24431, w24432, w24433, w24434, w24435, w24436, w24437, w24438, w24439, w24440, w24441, w24442, w24443, w24444, w24445, w24446, w24447, w24448, w24449, w24450, w24451, w24452, w24453, w24454, w24455, w24456, w24457, w24458, w24459, w24460, w24461, w24462, w24463, w24464, w24465, w24466, w24467, w24468, w24469, w24470, w24471, w24472, w24473, w24474, w24475, w24476, w24477, w24478, w24479, w24480, w24481, w24482, w24483, w24484, w24485, w24486, w24487, w24488, w24489, w24490, w24491, w24492, w24493, w24494, w24495, w24496, w24497, w24498, w24499, w24500, w24501, w24502, w24503, w24504, w24505, w24506, w24507, w24508, w24509, w24510, w24511, w24512, w24513, w24514, w24515, w24516, w24517, w24518, w24519, w24520, w24521, w24522, w24523, w24524, w24525, w24526, w24527, w24528, w24529, w24530, w24531, w24532, w24533, w24534, w24535, w24536, w24537, w24538, w24539, w24540, w24541, w24542, w24543, w24544, w24545, w24546, w24547, w24548, w24549, w24550, w24551, w24552, w24553, w24554, w24555, w24556, w24557, w24558, w24559, w24560, w24561, w24562, w24563, w24564, w24565, w24566, w24567, w24568, w24569, w24570, w24571, w24572, w24573, w24574, w24575, w24576, w24577, w24578, w24579, w24580, w24581, w24582, w24583, w24584, w24585, w24586, w24587, w24588, w24589, w24590, w24591, w24592, w24593, w24594, w24595, w24596, w24597, w24598, w24599, w24600, w24601, w24602, w24603, w24604, w24605, w24606, w24607, w24608, w24609, w24610, w24611, w24612, w24613, w24614, w24615, w24616, w24617, w24618, w24619, w24620, w24621, w24622, w24623, w24624, w24625, w24626, w24627, w24628, w24629, w24630, w24631, w24632, w24633, w24634, w24635, w24636, w24637, w24638, w24639, w24640, w24641, w24642, w24643, w24644, w24645, w24646, w24647, w24648, w24649, w24650, w24651, w24652, w24653, w24654, w24655, w24656, w24657, w24658, w24659, w24660, w24661, w24662, w24663, w24664, w24665, w24666, w24667, w24668, w24669, w24670, w24671, w24672, w24673, w24674, w24675, w24676, w24677, w24678, w24679, w24680, w24681, w24682, w24683, w24684, w24685, w24686, w24687, w24688, w24689, w24690, w24691, w24692, w24693, w24694, w24695, w24696, w24697, w24698, w24699, w24700, w24701, w24702, w24703, w24704, w24705, w24706, w24707, w24708, w24709, w24710, w24711, w24712, w24713, w24714, w24715, w24716, w24717, w24718, w24719, w24720, w24721, w24722, w24723, w24724, w24725, w24726, w24727, w24728, w24729, w24730, w24731, w24732, w24733, w24734, w24735, w24736, w24737, w24738, w24739, w24740, w24741, w24742, w24743, w24744, w24745, w24746, w24747, w24748, w24749, w24750, w24751, w24752, w24753, w24754, w24755, w24756, w24757, w24758, w24759, w24760, w24761, w24762, w24763, w24764, w24765, w24766, w24767, w24768, w24769, w24770, w24771, w24772, w24773, w24774, w24775, w24776, w24777, w24778, w24779, w24780, w24781, w24782, w24783, w24784, w24785, w24786, w24787, w24788, w24789, w24790, w24791, w24792, w24793, w24794, w24795, w24796, w24797, w24798, w24799, w24800, w24801, w24802, w24803, w24804, w24805, w24806, w24807, w24808, w24809, w24810, w24811, w24812, w24813, w24814, w24815, w24816, w24817, w24818, w24819, w24820, w24821, w24822, w24823, w24824, w24825, w24826, w24827, w24828, w24829, w24830, w24831, w24832, w24833, w24834, w24835, w24836, w24837, w24838, w24839, w24840, w24841, w24842, w24843, w24844, w24845, w24846, w24847, w24848, w24849, w24850, w24851, w24852, w24853, w24854, w24855, w24856, w24857, w24858, w24859, w24860, w24861, w24862, w24863, w24864, w24865, w24866, w24867, w24868, w24869, w24870, w24871, w24872, w24873, w24874, w24875, w24876, w24877, w24878, w24879, w24880, w24881, w24882, w24883, w24884, w24885, w24886, w24887, w24888, w24889, w24890, w24891, w24892, w24893, w24894, w24895, w24896, w24897, w24898, w24899, w24900, w24901, w24902, w24903, w24904, w24905, w24906, w24907, w24908, w24909, w24910, w24911, w24912, w24913, w24914, w24915, w24916, w24917, w24918, w24919, w24920, w24921, w24922, w24923, w24924, w24925, w24926, w24927, w24928, w24929, w24930, w24931, w24932, w24933, w24934, w24935, w24936, w24937, w24938, w24939, w24940, w24941, w24942, w24943, w24944, w24945, w24946, w24947, w24948, w24949, w24950, w24951, w24952, w24953, w24954, w24955, w24956, w24957, w24958, w24959, w24960, w24961, w24962, w24963, w24964, w24965, w24966, w24967, w24968, w24969, w24970, w24971, w24972, w24973, w24974, w24975, w24976, w24977, w24978, w24979, w24980, w24981, w24982, w24983, w24984, w24985, w24986, w24987, w24988, w24989, w24990, w24991, w24992, w24993, w24994, w24995, w24996, w24997, w24998, w24999, w25000, w25001, w25002, w25003, w25004, w25005, w25006, w25007, w25008, w25009, w25010, w25011, w25012, w25013, w25014, w25015, w25016, w25017, w25018, w25019, w25020, w25021, w25022, w25023, w25024, w25025, w25026, w25027, w25028, w25029, w25030, w25031, w25032, w25033, w25034, w25035, w25036, w25037, w25038, w25039, w25040, w25041, w25042, w25043, w25044, w25045, w25046, w25047, w25048, w25049, w25050, w25051, w25052, w25053, w25054, w25055, w25056, w25057, w25058, w25059, w25060, w25061, w25062, w25063, w25064, w25065, w25066, w25067, w25068, w25069, w25070, w25071, w25072, w25073, w25074, w25075, w25076, w25077, w25078, w25079, w25080, w25081, w25082, w25083, w25084, w25085, w25086, w25087, w25088, w25089, w25090, w25091, w25092, w25093, w25094, w25095, w25096, w25097, w25098, w25099, w25100, w25101, w25102, w25103, w25104, w25105, w25106, w25107, w25108, w25109, w25110, w25111, w25112, w25113, w25114, w25115, w25116, w25117, w25118, w25119, w25120, w25121, w25122, w25123, w25124, w25125, w25126, w25127, w25128, w25129, w25130, w25131, w25132, w25133, w25134, w25135, w25136, w25137, w25138, w25139, w25140, w25141, w25142, w25143, w25144, w25145, w25146, w25147, w25148, w25149, w25150, w25151, w25152, w25153, w25154, w25155, w25156, w25157, w25158, w25159, w25160, w25161, w25162, w25163, w25164, w25165, w25166, w25167, w25168, w25169, w25170, w25171, w25172, w25173, w25174, w25175, w25176, w25177, w25178, w25179, w25180, w25181, w25182, w25183, w25184, w25185, w25186, w25187, w25188, w25189, w25190, w25191, w25192, w25193, w25194, w25195, w25196, w25197, w25198, w25199, w25200, w25201, w25202, w25203, w25204, w25205, w25206, w25207, w25208, w25209, w25210, w25211, w25212, w25213, w25214, w25215, w25216, w25217, w25218, w25219, w25220, w25221, w25222, w25223, w25224, w25225, w25226, w25227, w25228, w25229, w25230, w25231, w25232, w25233, w25234, w25235, w25236, w25237, w25238, w25239, w25240, w25241, w25242, w25243, w25244, w25245, w25246, w25247, w25248, w25249, w25250, w25251, w25252, w25253, w25254, w25255, w25256, w25257, w25258, w25259, w25260, w25261, w25262, w25263, w25264, w25265, w25266, w25267, w25268, w25269, w25270, w25271, w25272, w25273, w25274, w25275, w25276, w25277, w25278, w25279, w25280, w25281, w25282, w25283, w25284, w25285, w25286, w25287, w25288, w25289, w25290, w25291, w25292, w25293, w25294, w25295, w25296, w25297, w25298, w25299, w25300, w25301, w25302, w25303, w25304, w25305, w25306, w25307, w25308, w25309, w25310, w25311, w25312, w25313, w25314, w25315, w25316, w25317, w25318, w25319, w25320, w25321, w25322, w25323, w25324, w25325, w25326, w25327, w25328, w25329, w25330, w25331, w25332, w25333, w25334, w25335, w25336, w25337, w25338, w25339, w25340, w25341, w25342, w25343, w25344, w25345, w25346, w25347, w25348, w25349, w25350, w25351, w25352, w25353, w25354, w25355, w25356, w25357, w25358, w25359, w25360, w25361, w25362, w25363, w25364, w25365, w25366, w25367, w25368, w25369, w25370, w25371, w25372, w25373, w25374, w25375, w25376, w25377, w25378, w25379, w25380, w25381, w25382, w25383, w25384, w25385, w25386, w25387, w25388, w25389, w25390, w25391, w25392, w25393, w25394, w25395, w25396, w25397, w25398, w25399, w25400, w25401, w25402, w25403, w25404, w25405, w25406, w25407, w25408, w25409, w25410, w25411, w25412, w25413, w25414, w25415, w25416, w25417, w25418, w25419, w25420, w25421, w25422, w25423, w25424, w25425, w25426, w25427, w25428, w25429, w25430, w25431, w25432, w25433, w25434, w25435, w25436, w25437, w25438, w25439, w25440, w25441, w25442, w25443, w25444, w25445, w25446, w25447, w25448, w25449, w25450, w25451, w25452, w25453, w25454, w25455, w25456, w25457, w25458, w25459, w25460, w25461, w25462, w25463, w25464, w25465, w25466, w25467, w25468, w25469, w25470, w25471, w25472, w25473, w25474, w25475, w25476, w25477, w25478, w25479, w25480, w25481, w25482, w25483, w25484, w25485, w25486, w25487, w25488, w25489, w25490, w25491, w25492, w25493, w25494, w25495, w25496, w25497, w25498, w25499, w25500, w25501, w25502, w25503, w25504, w25505, w25506, w25507, w25508, w25509, w25510, w25511, w25512, w25513, w25514, w25515, w25516, w25517, w25518, w25519, w25520, w25521, w25522, w25523, w25524, w25525, w25526, w25527, w25528, w25529, w25530, w25531, w25532, w25533, w25534, w25535, w25536, w25537, w25538, w25539, w25540, w25541, w25542, w25543, w25544, w25545, w25546, w25547, w25548, w25549, w25550, w25551, w25552, w25553, w25554, w25555, w25556, w25557, w25558, w25559, w25560, w25561, w25562, w25563, w25564, w25565, w25566, w25567, w25568, w25569, w25570, w25571, w25572, w25573, w25574, w25575, w25576, w25577, w25578, w25579, w25580, w25581, w25582, w25583, w25584, w25585, w25586, w25587, w25588, w25589, w25590, w25591, w25592, w25593, w25594, w25595, w25596, w25597, w25598, w25599, w25600, w25601, w25602, w25603, w25604, w25605, w25606, w25607, w25608, w25609, w25610, w25611, w25612, w25613, w25614, w25615, w25616, w25617, w25618, w25619, w25620, w25621, w25622, w25623, w25624, w25625, w25626, w25627, w25628, w25629, w25630, w25631, w25632, w25633, w25634, w25635, w25636, w25637, w25638, w25639, w25640, w25641, w25642, w25643, w25644, w25645, w25646, w25647, w25648, w25649, w25650, w25651, w25652, w25653, w25654, w25655, w25656, w25657, w25658, w25659, w25660, w25661, w25662, w25663, w25664, w25665, w25666, w25667, w25668, w25669, w25670, w25671, w25672, w25673, w25674, w25675, w25676, w25677, w25678, w25679, w25680, w25681, w25682, w25683, w25684, w25685, w25686, w25687, w25688, w25689, w25690, w25691, w25692, w25693, w25694, w25695, w25696, w25697, w25698, w25699, w25700, w25701, w25702, w25703, w25704, w25705, w25706, w25707, w25708, w25709, w25710, w25711, w25712, w25713, w25714, w25715, w25716, w25717, w25718, w25719, w25720, w25721, w25722, w25723, w25724, w25725, w25726, w25727, w25728, w25729, w25730, w25731, w25732, w25733, w25734, w25735, w25736, w25737, w25738, w25739, w25740, w25741, w25742, w25743, w25744, w25745, w25746, w25747, w25748, w25749, w25750, w25751, w25752, w25753, w25754, w25755, w25756, w25757, w25758, w25759, w25760, w25761, w25762, w25763, w25764, w25765, w25766, w25767, w25768, w25769, w25770, w25771, w25772, w25773, w25774, w25775, w25776, w25777, w25778, w25779, w25780, w25781, w25782, w25783, w25784, w25785, w25786, w25787, w25788, w25789, w25790, w25791, w25792, w25793, w25794, w25795, w25796, w25797, w25798, w25799, w25800, w25801, w25802, w25803, w25804, w25805, w25806, w25807, w25808, w25809, w25810, w25811, w25812, w25813, w25814, w25815, w25816, w25817, w25818, w25819, w25820, w25821, w25822, w25823, w25824, w25825, w25826, w25827, w25828, w25829, w25830, w25831, w25832, w25833, w25834, w25835, w25836, w25837, w25838, w25839, w25840, w25841, w25842, w25843, w25844, w25845, w25846, w25847, w25848, w25849, w25850, w25851, w25852, w25853, w25854, w25855, w25856, w25857, w25858, w25859, w25860, w25861, w25862, w25863, w25864, w25865, w25866, w25867, w25868, w25869, w25870, w25871, w25872, w25873, w25874, w25875, w25876, w25877, w25878, w25879, w25880, w25881, w25882, w25883, w25884, w25885, w25886, w25887, w25888, w25889, w25890, w25891, w25892, w25893, w25894, w25895, w25896, w25897, w25898, w25899, w25900, w25901, w25902, w25903, w25904, w25905, w25906, w25907, w25908, w25909, w25910, w25911, w25912, w25913, w25914, w25915, w25916, w25917, w25918, w25919, w25920, w25921, w25922, w25923, w25924, w25925, w25926, w25927, w25928, w25929, w25930, w25931, w25932, w25933, w25934, w25935, w25936, w25937, w25938, w25939, w25940, w25941, w25942, w25943, w25944, w25945, w25946, w25947, w25948, w25949, w25950, w25951, w25952, w25953, w25954, w25955, w25956, w25957, w25958, w25959, w25960, w25961, w25962, w25963, w25964, w25965, w25966, w25967, w25968, w25969, w25970, w25971, w25972, w25973, w25974, w25975, w25976, w25977, w25978, w25979, w25980, w25981, w25982, w25983, w25984, w25985, w25986, w25987, w25988, w25989, w25990, w25991, w25992, w25993, w25994, w25995, w25996, w25997, w25998, w25999, w26000, w26001, w26002, w26003, w26004, w26005, w26006, w26007, w26008, w26009, w26010, w26011, w26012, w26013, w26014, w26015, w26016, w26017, w26018, w26019, w26020, w26021, w26022, w26023, w26024, w26025, w26026, w26027, w26028, w26029, w26030, w26031, w26032, w26033, w26034, w26035, w26036, w26037, w26038, w26039, w26040, w26041, w26042, w26043, w26044, w26045, w26046, w26047, w26048, w26049, w26050, w26051, w26052, w26053, w26054, w26055, w26056, w26057, w26058, w26059, w26060, w26061, w26062, w26063, w26064, w26065, w26066, w26067, w26068, w26069, w26070, w26071, w26072, w26073, w26074, w26075, w26076, w26077, w26078, w26079, w26080, w26081, w26082, w26083, w26084, w26085, w26086, w26087, w26088, w26089, w26090, w26091, w26092, w26093, w26094, w26095, w26096, w26097, w26098, w26099, w26100, w26101, w26102, w26103, w26104, w26105, w26106, w26107, w26108, w26109, w26110, w26111, w26112, w26113, w26114, w26115, w26116, w26117, w26118, w26119, w26120, w26121, w26122, w26123, w26124, w26125, w26126, w26127, w26128, w26129, w26130, w26131, w26132, w26133, w26134, w26135, w26136, w26137, w26138, w26139, w26140, w26141, w26142, w26143, w26144, w26145, w26146, w26147, w26148, w26149, w26150, w26151, w26152, w26153, w26154, w26155, w26156, w26157, w26158, w26159, w26160, w26161, w26162, w26163, w26164, w26165, w26166, w26167, w26168, w26169, w26170, w26171, w26172, w26173, w26174, w26175, w26176, w26177, w26178, w26179, w26180, w26181, w26182, w26183, w26184, w26185, w26186, w26187, w26188, w26189, w26190, w26191, w26192, w26193, w26194, w26195, w26196, w26197, w26198, w26199, w26200, w26201, w26202, w26203, w26204, w26205, w26206, w26207, w26208, w26209, w26210, w26211, w26212, w26213, w26214, w26215, w26216, w26217, w26218, w26219, w26220, w26221, w26222, w26223, w26224, w26225, w26226, w26227, w26228, w26229, w26230, w26231, w26232, w26233, w26234, w26235, w26236, w26237, w26238, w26239, w26240, w26241, w26242, w26243, w26244, w26245, w26246, w26247, w26248, w26249, w26250, w26251, w26252, w26253, w26254, w26255, w26256, w26257, w26258, w26259, w26260, w26261, w26262, w26263, w26264, w26265, w26266, w26267, w26268, w26269, w26270, w26271, w26272, w26273, w26274, w26275, w26276, w26277, w26278, w26279, w26280, w26281, w26282, w26283, w26284, w26285, w26286, w26287, w26288, w26289, w26290, w26291, w26292, w26293, w26294, w26295, w26296, w26297, w26298, w26299, w26300, w26301, w26302, w26303, w26304, w26305, w26306, w26307, w26308, w26309, w26310, w26311, w26312, w26313, w26314, w26315, w26316, w26317, w26318, w26319, w26320, w26321, w26322, w26323, w26324, w26325, w26326, w26327, w26328, w26329, w26330, w26331, w26332, w26333, w26334, w26335, w26336, w26337, w26338, w26339, w26340, w26341, w26342, w26343, w26344, w26345, w26346, w26347, w26348, w26349, w26350, w26351, w26352, w26353, w26354, w26355, w26356, w26357, w26358, w26359, w26360, w26361, w26362, w26363, w26364, w26365, w26366, w26367, w26368, w26369, w26370, w26371, w26372, w26373, w26374, w26375, w26376, w26377, w26378, w26379, w26380, w26381, w26382, w26383, w26384, w26385, w26386, w26387, w26388, w26389, w26390, w26391, w26392, w26393, w26394, w26395, w26396, w26397, w26398, w26399, w26400, w26401, w26402, w26403, w26404, w26405, w26406, w26407, w26408, w26409, w26410, w26411, w26412, w26413, w26414, w26415, w26416, w26417, w26418, w26419, w26420, w26421, w26422, w26423, w26424, w26425, w26426, w26427, w26428, w26429, w26430, w26431, w26432, w26433, w26434, w26435, w26436, w26437, w26438, w26439, w26440, w26441, w26442, w26443, w26444, w26445, w26446, w26447, w26448, w26449, w26450, w26451, w26452, w26453, w26454, w26455, w26456, w26457, w26458, w26459, w26460, w26461, w26462, w26463, w26464, w26465, w26466, w26467, w26468, w26469, w26470, w26471, w26472, w26473, w26474, w26475, w26476, w26477, w26478, w26479, w26480, w26481, w26482, w26483, w26484, w26485, w26486, w26487, w26488, w26489, w26490, w26491, w26492, w26493, w26494, w26495, w26496, w26497, w26498, w26499, w26500, w26501, w26502, w26503, w26504, w26505, w26506, w26507, w26508, w26509, w26510, w26511, w26512, w26513, w26514, w26515, w26516, w26517, w26518, w26519, w26520, w26521, w26522, w26523, w26524, w26525, w26526, w26527, w26528, w26529, w26530, w26531, w26532, w26533, w26534, w26535, w26536, w26537, w26538, w26539, w26540, w26541, w26542, w26543, w26544, w26545, w26546, w26547, w26548, w26549, w26550, w26551, w26552, w26553, w26554, w26555, w26556, w26557, w26558, w26559, w26560, w26561, w26562, w26563, w26564, w26565, w26566, w26567, w26568, w26569, w26570, w26571, w26572, w26573, w26574, w26575, w26576, w26577, w26578, w26579, w26580, w26581, w26582, w26583, w26584, w26585, w26586, w26587, w26588, w26589, w26590, w26591, w26592, w26593, w26594, w26595, w26596, w26597, w26598, w26599, w26600, w26601, w26602, w26603, w26604, w26605, w26606, w26607, w26608, w26609, w26610, w26611, w26612, w26613, w26614, w26615, w26616, w26617, w26618, w26619, w26620, w26621, w26622, w26623, w26624, w26625, w26626, w26627, w26628, w26629, w26630, w26631, w26632, w26633, w26634, w26635, w26636, w26637, w26638, w26639, w26640, w26641, w26642, w26643, w26644, w26645, w26646, w26647, w26648, w26649, w26650, w26651, w26652, w26653, w26654, w26655, w26656, w26657, w26658, w26659, w26660, w26661, w26662, w26663, w26664, w26665, w26666, w26667, w26668, w26669, w26670, w26671, w26672, w26673, w26674, w26675, w26676, w26677, w26678, w26679, w26680, w26681, w26682, w26683, w26684, w26685, w26686, w26687, w26688, w26689, w26690, w26691, w26692, w26693, w26694, w26695, w26696, w26697, w26698, w26699, w26700, w26701, w26702, w26703, w26704, w26705, w26706, w26707, w26708, w26709, w26710, w26711, w26712, w26713, w26714, w26715, w26716, w26717, w26718, w26719, w26720, w26721, w26722, w26723, w26724, w26725, w26726, w26727, w26728, w26729, w26730, w26731, w26732, w26733, w26734, w26735, w26736, w26737, w26738, w26739, w26740, w26741, w26742, w26743, w26744, w26745, w26746, w26747, w26748, w26749, w26750, w26751, w26752, w26753, w26754, w26755, w26756, w26757, w26758, w26759, w26760, w26761, w26762, w26763, w26764, w26765, w26766, w26767, w26768, w26769, w26770, w26771, w26772, w26773, w26774, w26775, w26776, w26777, w26778, w26779, w26780, w26781, w26782, w26783, w26784, w26785, w26786, w26787, w26788, w26789, w26790, w26791, w26792, w26793, w26794, w26795, w26796, w26797, w26798, w26799, w26800, w26801, w26802, w26803, w26804, w26805, w26806, w26807, w26808, w26809, w26810, w26811, w26812, w26813, w26814, w26815, w26816, w26817, w26818, w26819, w26820, w26821, w26822, w26823, w26824, w26825, w26826, w26827, w26828, w26829, w26830, w26831, w26832, w26833, w26834, w26835, w26836, w26837, w26838, w26839, w26840, w26841, w26842, w26843, w26844, w26845, w26846, w26847, w26848, w26849, w26850, w26851, w26852, w26853, w26854, w26855, w26856, w26857, w26858, w26859, w26860, w26861, w26862, w26863, w26864, w26865, w26866, w26867, w26868, w26869, w26870, w26871, w26872, w26873, w26874, w26875, w26876, w26877, w26878, w26879, w26880, w26881, w26882, w26883, w26884, w26885, w26886, w26887, w26888, w26889, w26890, w26891, w26892, w26893, w26894, w26895, w26896, w26897, w26898, w26899, w26900, w26901, w26902, w26903, w26904, w26905, w26906, w26907, w26908, w26909, w26910, w26911, w26912, w26913, w26914, w26915, w26916, w26917, w26918, w26919, w26920, w26921, w26922, w26923, w26924, w26925, w26926, w26927, w26928, w26929, w26930, w26931, w26932, w26933, w26934, w26935, w26936, w26937, w26938, w26939, w26940, w26941, w26942, w26943, w26944, w26945, w26946, w26947, w26948, w26949, w26950, w26951, w26952, w26953, w26954, w26955, w26956, w26957, w26958, w26959, w26960, w26961, w26962, w26963, w26964, w26965, w26966, w26967, w26968, w26969, w26970, w26971, w26972, w26973, w26974, w26975, w26976, w26977, w26978, w26979, w26980, w26981, w26982, w26983, w26984, w26985, w26986, w26987, w26988, w26989, w26990, w26991, w26992, w26993, w26994, w26995, w26996, w26997, w26998, w26999, w27000, w27001, w27002, w27003, w27004, w27005, w27006, w27007, w27008, w27009, w27010, w27011, w27012, w27013, w27014, w27015, w27016, w27017, w27018, w27019, w27020, w27021, w27022, w27023, w27024, w27025, w27026, w27027, w27028, w27029, w27030, w27031, w27032, w27033, w27034, w27035, w27036, w27037, w27038, w27039, w27040, w27041, w27042, w27043, w27044, w27045, w27046, w27047, w27048, w27049, w27050, w27051, w27052, w27053, w27054, w27055, w27056, w27057, w27058, w27059, w27060, w27061, w27062, w27063, w27064, w27065, w27066, w27067, w27068, w27069, w27070, w27071, w27072, w27073, w27074, w27075, w27076, w27077, w27078, w27079, w27080, w27081, w27082, w27083, w27084, w27085, w27086, w27087, w27088, w27089, w27090, w27091, w27092, w27093, w27094, w27095, w27096, w27097, w27098, w27099, w27100, w27101, w27102, w27103, w27104, w27105, w27106, w27107, w27108, w27109, w27110, w27111, w27112, w27113, w27114, w27115, w27116, w27117, w27118, w27119, w27120, w27121, w27122, w27123, w27124, w27125, w27126, w27127, w27128, w27129, w27130, w27131, w27132, w27133, w27134, w27135, w27136, w27137, w27138, w27139, w27140, w27141, w27142, w27143, w27144, w27145, w27146, w27147, w27148, w27149, w27150, w27151, w27152, w27153, w27154, w27155, w27156, w27157, w27158, w27159, w27160, w27161, w27162, w27163, w27164, w27165, w27166, w27167, w27168, w27169, w27170, w27171, w27172, w27173, w27174, w27175, w27176, w27177, w27178, w27179, w27180, w27181, w27182, w27183, w27184, w27185, w27186, w27187, w27188, w27189, w27190, w27191, w27192, w27193, w27194, w27195, w27196, w27197, w27198, w27199, w27200, w27201, w27202, w27203, w27204, w27205, w27206, w27207, w27208, w27209, w27210, w27211, w27212, w27213, w27214, w27215, w27216, w27217, w27218, w27219, w27220, w27221, w27222, w27223, w27224, w27225, w27226, w27227, w27228, w27229, w27230, w27231, w27232, w27233, w27234, w27235, w27236, w27237, w27238, w27239, w27240, w27241, w27242, w27243, w27244, w27245, w27246, w27247, w27248, w27249, w27250, w27251, w27252, w27253, w27254, w27255, w27256, w27257, w27258, w27259, w27260, w27261, w27262, w27263, w27264, w27265, w27266, w27267, w27268, w27269, w27270, w27271, w27272, w27273, w27274, w27275, w27276, w27277, w27278, w27279, w27280, w27281, w27282, w27283, w27284, w27285, w27286, w27287, w27288, w27289, w27290, w27291, w27292, w27293, w27294, w27295, w27296, w27297, w27298, w27299, w27300, w27301, w27302, w27303, w27304, w27305, w27306, w27307, w27308, w27309, w27310, w27311, w27312, w27313, w27314, w27315, w27316, w27317, w27318, w27319, w27320, w27321, w27322, w27323, w27324, w27325, w27326, w27327, w27328, w27329, w27330, w27331, w27332, w27333, w27334, w27335, w27336, w27337, w27338, w27339, w27340, w27341, w27342, w27343, w27344, w27345, w27346, w27347, w27348, w27349, w27350, w27351, w27352, w27353, w27354, w27355, w27356, w27357, w27358, w27359, w27360, w27361, w27362, w27363, w27364, w27365, w27366, w27367, w27368, w27369, w27370, w27371, w27372, w27373, w27374, w27375, w27376, w27377, w27378, w27379, w27380, w27381, w27382, w27383, w27384, w27385, w27386, w27387, w27388, w27389, w27390, w27391, w27392, w27393, w27394, w27395, w27396, w27397, w27398, w27399, w27400, w27401, w27402, w27403, w27404, w27405, w27406, w27407, w27408, w27409, w27410, w27411, w27412, w27413, w27414, w27415, w27416, w27417, w27418, w27419, w27420, w27421, w27422, w27423, w27424, w27425, w27426, w27427, w27428, w27429, w27430, w27431, w27432, w27433, w27434, w27435, w27436, w27437, w27438, w27439, w27440, w27441, w27442, w27443, w27444, w27445, w27446, w27447, w27448, w27449, w27450, w27451, w27452, w27453, w27454, w27455, w27456, w27457, w27458, w27459, w27460, w27461, w27462, w27463, w27464, w27465, w27466, w27467, w27468, w27469, w27470, w27471, w27472, w27473, w27474, w27475, w27476, w27477, w27478, w27479, w27480, w27481, w27482, w27483, w27484, w27485, w27486, w27487, w27488, w27489, w27490, w27491, w27492, w27493, w27494, w27495, w27496, w27497, w27498, w27499, w27500, w27501, w27502, w27503, w27504, w27505, w27506, w27507, w27508, w27509, w27510, w27511, w27512, w27513, w27514, w27515, w27516, w27517, w27518, w27519, w27520, w27521, w27522, w27523, w27524, w27525, w27526, w27527, w27528, w27529, w27530, w27531, w27532, w27533, w27534, w27535, w27536, w27537, w27538, w27539, w27540, w27541, w27542, w27543, w27544, w27545, w27546, w27547, w27548, w27549, w27550, w27551, w27552, w27553, w27554, w27555, w27556, w27557, w27558, w27559, w27560, w27561, w27562, w27563, w27564, w27565, w27566, w27567, w27568, w27569, w27570, w27571, w27572, w27573, w27574, w27575, w27576, w27577, w27578, w27579, w27580, w27581, w27582, w27583, w27584, w27585, w27586, w27587, w27588, w27589, w27590, w27591, w27592, w27593, w27594, w27595, w27596, w27597, w27598, w27599, w27600, w27601, w27602, w27603, w27604, w27605, w27606, w27607, w27608, w27609, w27610, w27611, w27612, w27613, w27614, w27615, w27616, w27617, w27618, w27619, w27620, w27621, w27622, w27623, w27624, w27625, w27626, w27627, w27628, w27629, w27630, w27631, w27632, w27633, w27634, w27635, w27636, w27637, w27638, w27639, w27640, w27641, w27642, w27643, w27644, w27645, w27646, w27647, w27648, w27649, w27650, w27651, w27652, w27653, w27654, w27655, w27656, w27657, w27658, w27659, w27660, w27661, w27662, w27663, w27664, w27665, w27666, w27667, w27668, w27669, w27670, w27671, w27672, w27673, w27674, w27675, w27676, w27677, w27678, w27679, w27680, w27681, w27682, w27683, w27684, w27685, w27686, w27687, w27688, w27689, w27690, w27691, w27692, w27693, w27694, w27695, w27696, w27697, w27698, w27699, w27700, w27701, w27702, w27703, w27704, w27705, w27706, w27707, w27708, w27709, w27710, w27711, w27712, w27713, w27714, w27715, w27716, w27717, w27718, w27719, w27720, w27721, w27722, w27723, w27724, w27725, w27726, w27727, w27728, w27729, w27730, w27731, w27732, w27733, w27734, w27735, w27736, w27737, w27738, w27739, w27740, w27741, w27742, w27743, w27744, w27745, w27746, w27747, w27748, w27749, w27750, w27751, w27752, w27753, w27754, w27755, w27756, w27757, w27758, w27759, w27760, w27761, w27762, w27763, w27764, w27765, w27766, w27767, w27768, w27769, w27770, w27771, w27772, w27773, w27774, w27775, w27776, w27777, w27778, w27779, w27780, w27781, w27782, w27783, w27784, w27785, w27786, w27787, w27788, w27789, w27790, w27791, w27792, w27793, w27794, w27795, w27796, w27797, w27798, w27799, w27800, w27801, w27802, w27803, w27804, w27805, w27806, w27807, w27808, w27809, w27810, w27811, w27812, w27813, w27814, w27815, w27816, w27817, w27818, w27819, w27820, w27821, w27822, w27823, w27824, w27825, w27826, w27827, w27828, w27829, w27830, w27831, w27832, w27833, w27834, w27835, w27836, w27837, w27838, w27839, w27840, w27841, w27842, w27843, w27844, w27845, w27846, w27847, w27848, w27849, w27850, w27851, w27852, w27853, w27854, w27855, w27856, w27857, w27858, w27859, w27860, w27861, w27862, w27863, w27864, w27865, w27866, w27867, w27868, w27869, w27870, w27871, w27872, w27873, w27874, w27875, w27876, w27877, w27878, w27879, w27880, w27881, w27882, w27883, w27884, w27885, w27886, w27887, w27888, w27889, w27890, w27891, w27892, w27893, w27894, w27895, w27896, w27897, w27898, w27899, w27900, w27901, w27902, w27903, w27904, w27905, w27906, w27907, w27908, w27909, w27910, w27911, w27912, w27913, w27914, w27915, w27916, w27917, w27918, w27919, w27920, w27921, w27922, w27923, w27924, w27925, w27926, w27927, w27928, w27929, w27930, w27931, w27932, w27933, w27934, w27935, w27936, w27937, w27938, w27939, w27940, w27941, w27942, w27943, w27944, w27945, w27946, w27947, w27948, w27949, w27950, w27951, w27952, w27953, w27954, w27955, w27956, w27957, w27958, w27959, w27960, w27961, w27962, w27963, w27964, w27965, w27966, w27967, w27968, w27969, w27970, w27971, w27972, w27973, w27974, w27975, w27976, w27977, w27978, w27979, w27980, w27981, w27982, w27983, w27984, w27985, w27986, w27987, w27988, w27989, w27990, w27991, w27992, w27993, w27994, w27995, w27996, w27997, w27998, w27999, w28000, w28001, w28002, w28003, w28004, w28005, w28006, w28007, w28008, w28009, w28010, w28011, w28012, w28013, w28014, w28015, w28016, w28017, w28018, w28019, w28020, w28021, w28022, w28023, w28024, w28025, w28026, w28027, w28028, w28029, w28030, w28031, w28032, w28033, w28034, w28035, w28036, w28037, w28038, w28039, w28040, w28041, w28042, w28043, w28044, w28045, w28046, w28047, w28048, w28049, w28050, w28051, w28052, w28053, w28054, w28055, w28056, w28057, w28058, w28059, w28060, w28061, w28062, w28063, w28064, w28065, w28066, w28067, w28068, w28069, w28070, w28071, w28072, w28073, w28074, w28075, w28076, w28077, w28078, w28079, w28080, w28081, w28082, w28083, w28084, w28085, w28086, w28087, w28088, w28089, w28090, w28091, w28092, w28093, w28094, w28095, w28096, w28097, w28098, w28099, w28100, w28101, w28102, w28103, w28104, w28105, w28106, w28107, w28108, w28109, w28110, w28111, w28112, w28113, w28114, w28115, w28116, w28117, w28118, w28119, w28120, w28121, w28122, w28123, w28124, w28125, w28126, w28127, w28128, w28129, w28130, w28131, w28132, w28133, w28134, w28135, w28136, w28137, w28138, w28139, w28140, w28141, w28142, w28143, w28144, w28145, w28146, w28147, w28148, w28149, w28150, w28151, w28152, w28153, w28154, w28155, w28156, w28157, w28158, w28159, w28160, w28161, w28162, w28163, w28164, w28165, w28166, w28167, w28168, w28169, w28170, w28171, w28172, w28173, w28174, w28175, w28176, w28177, w28178, w28179, w28180, w28181, w28182, w28183, w28184, w28185, w28186, w28187, w28188, w28189, w28190, w28191, w28192, w28193, w28194, w28195, w28196, w28197, w28198, w28199, w28200, w28201, w28202, w28203, w28204, w28205, w28206, w28207, w28208, w28209, w28210, w28211, w28212, w28213, w28214, w28215, w28216, w28217, w28218, w28219, w28220, w28221, w28222, w28223, w28224, w28225, w28226, w28227, w28228, w28229, w28230, w28231, w28232, w28233, w28234, w28235, w28236, w28237, w28238, w28239, w28240, w28241, w28242, w28243, w28244, w28245, w28246, w28247, w28248, w28249, w28250, w28251, w28252, w28253, w28254, w28255, w28256, w28257, w28258, w28259, w28260, w28261, w28262, w28263, w28264, w28265, w28266, w28267, w28268, w28269, w28270, w28271, w28272, w28273, w28274, w28275, w28276, w28277, w28278, w28279, w28280, w28281, w28282, w28283, w28284, w28285, w28286, w28287, w28288, w28289, w28290, w28291, w28292, w28293, w28294, w28295, w28296, w28297, w28298, w28299, w28300, w28301, w28302, w28303, w28304, w28305, w28306, w28307, w28308, w28309, w28310, w28311, w28312, w28313, w28314, w28315, w28316, w28317, w28318, w28319, w28320, w28321, w28322, w28323, w28324, w28325, w28326, w28327, w28328, w28329, w28330, w28331, w28332, w28333, w28334, w28335, w28336, w28337, w28338, w28339, w28340, w28341, w28342, w28343, w28344, w28345, w28346, w28347, w28348, w28349, w28350, w28351, w28352, w28353, w28354, w28355, w28356, w28357, w28358, w28359, w28360, w28361, w28362, w28363, w28364, w28365, w28366, w28367, w28368, w28369, w28370, w28371, w28372, w28373, w28374, w28375, w28376, w28377, w28378, w28379, w28380, w28381, w28382, w28383, w28384, w28385, w28386, w28387, w28388, w28389, w28390, w28391, w28392, w28393, w28394, w28395, w28396, w28397, w28398, w28399, w28400, w28401, w28402, w28403, w28404, w28405, w28406, w28407, w28408, w28409, w28410, w28411, w28412, w28413, w28414, w28415, w28416, w28417, w28418, w28419, w28420, w28421, w28422, w28423, w28424, w28425, w28426, w28427, w28428, w28429, w28430, w28431, w28432, w28433, w28434, w28435, w28436, w28437, w28438, w28439, w28440, w28441, w28442, w28443, w28444, w28445, w28446, w28447, w28448, w28449, w28450, w28451, w28452, w28453, w28454, w28455, w28456, w28457, w28458, w28459, w28460, w28461, w28462, w28463, w28464, w28465, w28466, w28467, w28468, w28469, w28470, w28471, w28472, w28473, w28474, w28475, w28476, w28477, w28478, w28479, w28480, w28481, w28482, w28483, w28484, w28485, w28486, w28487, w28488, w28489, w28490, w28491, w28492, w28493, w28494, w28495, w28496, w28497, w28498, w28499, w28500, w28501, w28502, w28503, w28504, w28505, w28506, w28507, w28508, w28509, w28510, w28511, w28512, w28513, w28514, w28515, w28516, w28517, w28518, w28519, w28520, w28521, w28522, w28523, w28524, w28525, w28526, w28527, w28528, w28529, w28530, w28531, w28532, w28533, w28534, w28535, w28536, w28537, w28538, w28539, w28540, w28541, w28542, w28543, w28544, w28545, w28546, w28547, w28548, w28549, w28550, w28551, w28552, w28553, w28554, w28555, w28556, w28557, w28558, w28559, w28560, w28561, w28562, w28563, w28564, w28565, w28566, w28567, w28568, w28569, w28570, w28571, w28572, w28573, w28574, w28575, w28576, w28577, w28578, w28579, w28580, w28581, w28582, w28583, w28584, w28585, w28586, w28587, w28588, w28589, w28590, w28591, w28592, w28593, w28594, w28595, w28596, w28597, w28598, w28599, w28600, w28601, w28602, w28603, w28604, w28605, w28606, w28607, w28608, w28609, w28610, w28611, w28612, w28613, w28614, w28615, w28616, w28617, w28618, w28619, w28620, w28621, w28622, w28623, w28624, w28625, w28626, w28627, w28628, w28629, w28630, w28631, w28632, w28633, w28634, w28635, w28636, w28637, w28638, w28639, w28640, w28641, w28642, w28643, w28644, w28645, w28646, w28647, w28648, w28649, w28650, w28651, w28652, w28653, w28654, w28655, w28656, w28657, w28658, w28659, w28660, w28661, w28662, w28663, w28664, w28665, w28666, w28667, w28668, w28669, w28670, w28671, w28672, w28673, w28674, w28675, w28676, w28677, w28678, w28679, w28680, w28681, w28682, w28683, w28684, w28685, w28686, w28687, w28688, w28689, w28690, w28691, w28692, w28693, w28694, w28695, w28696, w28697, w28698, w28699, w28700, w28701, w28702, w28703, w28704, w28705, w28706, w28707, w28708, w28709, w28710, w28711, w28712, w28713, w28714, w28715, w28716, w28717, w28718, w28719, w28720, w28721, w28722, w28723, w28724, w28725, w28726, w28727, w28728, w28729, w28730, w28731, w28732, w28733, w28734, w28735, w28736, w28737, w28738, w28739, w28740, w28741, w28742, w28743, w28744, w28745, w28746, w28747, w28748, w28749, w28750, w28751, w28752, w28753, w28754, w28755, w28756, w28757, w28758, w28759, w28760, w28761, w28762, w28763, w28764, w28765, w28766, w28767, w28768, w28769, w28770, w28771, w28772, w28773, w28774, w28775, w28776, w28777, w28778, w28779, w28780, w28781, w28782, w28783, w28784, w28785, w28786, w28787, w28788, w28789, w28790, w28791, w28792, w28793, w28794, w28795, w28796, w28797, w28798, w28799, w28800, w28801, w28802, w28803, w28804, w28805, w28806, w28807, w28808, w28809, w28810, w28811, w28812, w28813, w28814, w28815, w28816, w28817, w28818, w28819, w28820, w28821, w28822, w28823, w28824, w28825, w28826, w28827, w28828, w28829, w28830, w28831, w28832, w28833, w28834, w28835, w28836, w28837, w28838, w28839, w28840, w28841, w28842, w28843, w28844, w28845, w28846, w28847, w28848, w28849, w28850, w28851, w28852, w28853, w28854, w28855, w28856, w28857, w28858, w28859, w28860, w28861, w28862, w28863, w28864, w28865, w28866, w28867, w28868, w28869, w28870, w28871, w28872, w28873, w28874, w28875, w28876, w28877, w28878, w28879, w28880, w28881, w28882, w28883, w28884, w28885, w28886, w28887, w28888, w28889, w28890, w28891, w28892, w28893, w28894, w28895, w28896, w28897, w28898, w28899, w28900, w28901, w28902, w28903, w28904, w28905, w28906, w28907, w28908, w28909, w28910, w28911, w28912, w28913, w28914, w28915, w28916, w28917, w28918, w28919, w28920, w28921, w28922, w28923, w28924, w28925, w28926, w28927, w28928, w28929, w28930, w28931, w28932, w28933, w28934, w28935, w28936, w28937, w28938, w28939, w28940, w28941, w28942, w28943, w28944, w28945, w28946, w28947, w28948, w28949, w28950, w28951, w28952, w28953, w28954, w28955, w28956, w28957, w28958, w28959, w28960, w28961, w28962, w28963, w28964, w28965, w28966, w28967, w28968, w28969, w28970, w28971, w28972, w28973, w28974, w28975, w28976, w28977, w28978, w28979, w28980, w28981, w28982, w28983, w28984, w28985, w28986, w28987, w28988, w28989, w28990, w28991, w28992, w28993, w28994, w28995, w28996, w28997, w28998, w28999, w29000, w29001, w29002, w29003, w29004, w29005, w29006, w29007, w29008, w29009, w29010, w29011, w29012, w29013, w29014, w29015, w29016, w29017, w29018, w29019, w29020, w29021, w29022, w29023, w29024, w29025, w29026, w29027, w29028, w29029, w29030, w29031, w29032, w29033, w29034, w29035, w29036, w29037, w29038, w29039, w29040, w29041, w29042, w29043, w29044, w29045, w29046, w29047, w29048, w29049, w29050, w29051, w29052, w29053, w29054, w29055, w29056, w29057, w29058, w29059, w29060, w29061, w29062, w29063, w29064, w29065, w29066, w29067, w29068, w29069, w29070, w29071, w29072, w29073, w29074, w29075, w29076, w29077, w29078, w29079, w29080, w29081, w29082, w29083, w29084, w29085, w29086, w29087, w29088, w29089, w29090, w29091, w29092, w29093, w29094, w29095, w29096, w29097, w29098, w29099, w29100, w29101, w29102, w29103, w29104, w29105, w29106, w29107, w29108, w29109, w29110, w29111, w29112, w29113, w29114, w29115, w29116, w29117, w29118, w29119, w29120, w29121, w29122, w29123, w29124, w29125, w29126, w29127, w29128, w29129, w29130, w29131, w29132, w29133, w29134, w29135, w29136, w29137, w29138, w29139, w29140, w29141, w29142, w29143, w29144, w29145, w29146, w29147, w29148, w29149, w29150, w29151, w29152, w29153, w29154, w29155, w29156, w29157, w29158, w29159, w29160, w29161, w29162, w29163, w29164, w29165, w29166, w29167, w29168, w29169, w29170, w29171, w29172, w29173, w29174, w29175, w29176, w29177, w29178, w29179, w29180, w29181, w29182, w29183, w29184, w29185, w29186, w29187, w29188, w29189, w29190, w29191, w29192, w29193, w29194, w29195, w29196, w29197, w29198, w29199, w29200, w29201, w29202, w29203, w29204, w29205, w29206, w29207, w29208, w29209, w29210, w29211, w29212, w29213, w29214, w29215, w29216, w29217, w29218, w29219, w29220, w29221, w29222, w29223, w29224, w29225, w29226, w29227, w29228, w29229, w29230, w29231, w29232, w29233, w29234, w29235, w29236, w29237, w29238, w29239, w29240, w29241, w29242, w29243, w29244, w29245, w29246, w29247, w29248, w29249, w29250, w29251, w29252, w29253, w29254, w29255, w29256, w29257, w29258, w29259, w29260, w29261, w29262, w29263, w29264, w29265, w29266, w29267, w29268, w29269, w29270, w29271, w29272, w29273, w29274, w29275, w29276, w29277, w29278, w29279, w29280, w29281, w29282, w29283, w29284, w29285, w29286, w29287, w29288, w29289, w29290, w29291, w29292, w29293, w29294, w29295, w29296, w29297, w29298, w29299, w29300, w29301, w29302, w29303, w29304, w29305, w29306, w29307, w29308, w29309, w29310, w29311, w29312, w29313, w29314, w29315, w29316, w29317, w29318, w29319, w29320, w29321, w29322, w29323, w29324, w29325, w29326, w29327, w29328, w29329, w29330, w29331, w29332, w29333, w29334, w29335, w29336, w29337, w29338, w29339, w29340, w29341, w29342, w29343, w29344, w29345, w29346, w29347, w29348, w29349, w29350, w29351, w29352, w29353, w29354, w29355, w29356, w29357, w29358, w29359, w29360, w29361, w29362, w29363, w29364, w29365, w29366, w29367, w29368, w29369, w29370, w29371, w29372, w29373, w29374, w29375, w29376, w29377, w29378, w29379, w29380, w29381, w29382, w29383, w29384, w29385, w29386, w29387, w29388, w29389, w29390, w29391, w29392, w29393, w29394, w29395, w29396, w29397, w29398, w29399, w29400, w29401, w29402, w29403, w29404, w29405, w29406, w29407, w29408, w29409, w29410, w29411, w29412, w29413, w29414, w29415, w29416, w29417, w29418, w29419, w29420, w29421, w29422, w29423, w29424, w29425, w29426, w29427, w29428, w29429, w29430, w29431, w29432, w29433, w29434, w29435, w29436, w29437, w29438, w29439, w29440, w29441, w29442, w29443, w29444, w29445, w29446, w29447, w29448, w29449, w29450, w29451, w29452, w29453, w29454, w29455, w29456, w29457, w29458, w29459, w29460, w29461, w29462, w29463, w29464, w29465, w29466, w29467, w29468, w29469, w29470, w29471, w29472, w29473, w29474, w29475, w29476, w29477, w29478, w29479, w29480, w29481, w29482, w29483, w29484, w29485, w29486, w29487, w29488, w29489, w29490, w29491, w29492, w29493, w29494, w29495, w29496, w29497, w29498, w29499, w29500, w29501, w29502, w29503, w29504, w29505, w29506, w29507, w29508, w29509, w29510, w29511, w29512, w29513, w29514, w29515, w29516, w29517, w29518, w29519, w29520, w29521, w29522, w29523, w29524, w29525, w29526, w29527, w29528, w29529, w29530, w29531, w29532, w29533, w29534, w29535, w29536, w29537, w29538, w29539, w29540, w29541, w29542, w29543, w29544, w29545, w29546, w29547, w29548, w29549, w29550, w29551, w29552, w29553, w29554, w29555, w29556, w29557, w29558, w29559, w29560, w29561, w29562, w29563, w29564, w29565, w29566, w29567, w29568, w29569, w29570, w29571, w29572, w29573, w29574, w29575, w29576, w29577, w29578, w29579, w29580, w29581, w29582, w29583, w29584, w29585, w29586, w29587, w29588, w29589, w29590, w29591, w29592, w29593, w29594, w29595, w29596, w29597, w29598, w29599, w29600, w29601, w29602, w29603, w29604, w29605, w29606, w29607, w29608, w29609, w29610, w29611, w29612, w29613, w29614, w29615, w29616, w29617, w29618, w29619, w29620, w29621, w29622, w29623, w29624, w29625, w29626, w29627, w29628, w29629, w29630, w29631, w29632, w29633, w29634, w29635, w29636, w29637, w29638, w29639, w29640, w29641, w29642, w29643, w29644, w29645, w29646, w29647, w29648, w29649, w29650, w29651, w29652, w29653, w29654, w29655, w29656, w29657, w29658, w29659, w29660, w29661, w29662, w29663, w29664, w29665, w29666, w29667, w29668, w29669, w29670, w29671, w29672, w29673, w29674, w29675, w29676, w29677, w29678, w29679, w29680, w29681, w29682, w29683, w29684, w29685, w29686, w29687, w29688, w29689, w29690, w29691, w29692, w29693, w29694, w29695, w29696, w29697, w29698, w29699, w29700, w29701, w29702, w29703, w29704, w29705, w29706, w29707, w29708, w29709, w29710, w29711, w29712, w29713, w29714, w29715, w29716, w29717, w29718, w29719, w29720, w29721, w29722, w29723, w29724, w29725, w29726, w29727, w29728, w29729, w29730, w29731, w29732, w29733, w29734, w29735, w29736, w29737, w29738, w29739, w29740, w29741, w29742, w29743, w29744, w29745, w29746, w29747, w29748, w29749, w29750, w29751, w29752, w29753, w29754, w29755, w29756, w29757, w29758, w29759, w29760, w29761, w29762, w29763, w29764, w29765, w29766, w29767, w29768, w29769, w29770, w29771, w29772, w29773, w29774, w29775, w29776, w29777, w29778, w29779, w29780, w29781, w29782, w29783, w29784, w29785, w29786, w29787, w29788, w29789, w29790, w29791, w29792, w29793, w29794, w29795, w29796, w29797, w29798, w29799, w29800, w29801, w29802, w29803, w29804, w29805, w29806, w29807, w29808, w29809, w29810, w29811, w29812, w29813, w29814, w29815, w29816, w29817, w29818, w29819, w29820, w29821, w29822, w29823, w29824, w29825, w29826, w29827, w29828, w29829, w29830, w29831, w29832, w29833, w29834, w29835, w29836, w29837, w29838, w29839, w29840, w29841, w29842, w29843, w29844, w29845, w29846, w29847, w29848, w29849, w29850, w29851, w29852, w29853, w29854, w29855, w29856, w29857, w29858, w29859, w29860, w29861, w29862, w29863, w29864, w29865, w29866, w29867, w29868, w29869, w29870, w29871, w29872, w29873, w29874, w29875, w29876, w29877, w29878, w29879, w29880, w29881, w29882, w29883, w29884, w29885, w29886, w29887, w29888, w29889, w29890, w29891, w29892, w29893, w29894, w29895, w29896, w29897, w29898, w29899, w29900, w29901, w29902, w29903, w29904, w29905, w29906, w29907, w29908, w29909, w29910, w29911, w29912, w29913, w29914, w29915, w29916, w29917, w29918, w29919, w29920, w29921, w29922, w29923, w29924, w29925, w29926, w29927, w29928, w29929, w29930, w29931, w29932, w29933, w29934, w29935, w29936, w29937, w29938, w29939, w29940, w29941, w29942, w29943, w29944, w29945, w29946, w29947, w29948, w29949, w29950, w29951, w29952, w29953, w29954, w29955, w29956, w29957, w29958, w29959, w29960, w29961, w29962, w29963, w29964, w29965, w29966, w29967, w29968, w29969, w29970, w29971, w29972, w29973, w29974, w29975, w29976, w29977, w29978, w29979, w29980, w29981, w29982, w29983, w29984, w29985, w29986, w29987, w29988, w29989, w29990, w29991, w29992, w29993, w29994, w29995, w29996, w29997, w29998, w29999, w30000, w30001, w30002, w30003, w30004, w30005, w30006, w30007, w30008, w30009, w30010, w30011, w30012, w30013, w30014, w30015, w30016, w30017, w30018, w30019, w30020, w30021, w30022, w30023, w30024, w30025, w30026, w30027, w30028, w30029, w30030, w30031, w30032, w30033, w30034, w30035, w30036, w30037, w30038, w30039, w30040, w30041, w30042, w30043, w30044, w30045, w30046, w30047, w30048, w30049, w30050, w30051, w30052, w30053, w30054, w30055, w30056, w30057, w30058, w30059, w30060, w30061, w30062, w30063, w30064, w30065, w30066, w30067, w30068, w30069, w30070, w30071, w30072, w30073, w30074, w30075, w30076, w30077, w30078, w30079, w30080, w30081, w30082, w30083, w30084, w30085, w30086, w30087, w30088, w30089, w30090, w30091, w30092, w30093, w30094, w30095, w30096, w30097, w30098, w30099, w30100, w30101, w30102, w30103, w30104, w30105, w30106, w30107, w30108, w30109, w30110, w30111, w30112, w30113, w30114, w30115, w30116, w30117, w30118, w30119, w30120, w30121, w30122, w30123, w30124, w30125, w30126, w30127, w30128, w30129, w30130, w30131, w30132, w30133, w30134, w30135, w30136, w30137, w30138, w30139, w30140, w30141, w30142, w30143, w30144, w30145, w30146, w30147, w30148, w30149, w30150, w30151, w30152, w30153, w30154, w30155, w30156, w30157, w30158, w30159, w30160, w30161, w30162, w30163, w30164, w30165, w30166, w30167, w30168, w30169, w30170, w30171, w30172, w30173, w30174, w30175, w30176, w30177, w30178, w30179, w30180, w30181, w30182, w30183, w30184, w30185, w30186, w30187, w30188, w30189, w30190, w30191, w30192, w30193, w30194, w30195, w30196, w30197, w30198, w30199, w30200, w30201, w30202, w30203, w30204, w30205, w30206, w30207, w30208, w30209, w30210, w30211, w30212, w30213, w30214, w30215, w30216, w30217, w30218, w30219, w30220, w30221, w30222, w30223, w30224, w30225, w30226, w30227, w30228, w30229, w30230, w30231, w30232, w30233, w30234, w30235, w30236, w30237, w30238, w30239, w30240, w30241, w30242, w30243, w30244, w30245, w30246, w30247, w30248, w30249, w30250, w30251, w30252, w30253, w30254, w30255, w30256, w30257, w30258, w30259, w30260, w30261, w30262, w30263, w30264, w30265, w30266, w30267, w30268, w30269, w30270, w30271, w30272, w30273, w30274, w30275, w30276, w30277, w30278, w30279, w30280, w30281, w30282, w30283, w30284, w30285, w30286, w30287, w30288, w30289, w30290, w30291, w30292, w30293, w30294, w30295, w30296, w30297, w30298, w30299, w30300, w30301, w30302, w30303, w30304, w30305, w30306, w30307, w30308, w30309, w30310, w30311, w30312, w30313, w30314, w30315, w30316, w30317, w30318, w30319, w30320, w30321, w30322, w30323, w30324, w30325, w30326, w30327, w30328, w30329, w30330, w30331, w30332, w30333, w30334, w30335, w30336, w30337, w30338, w30339, w30340, w30341, w30342, w30343, w30344, w30345, w30346, w30347, w30348, w30349, w30350, w30351, w30352, w30353, w30354, w30355, w30356, w30357, w30358, w30359, w30360, w30361, w30362, w30363, w30364, w30365, w30366, w30367, w30368, w30369, w30370, w30371, w30372, w30373, w30374, w30375, w30376, w30377, w30378, w30379, w30380, w30381, w30382, w30383, w30384, w30385, w30386, w30387, w30388, w30389, w30390, w30391, w30392, w30393, w30394, w30395, w30396, w30397, w30398, w30399, w30400, w30401, w30402, w30403, w30404, w30405, w30406, w30407, w30408, w30409, w30410, w30411, w30412, w30413, w30414, w30415, w30416, w30417, w30418, w30419, w30420, w30421, w30422, w30423, w30424, w30425, w30426, w30427, w30428, w30429, w30430, w30431, w30432, w30433, w30434, w30435, w30436, w30437, w30438, w30439, w30440, w30441, w30442, w30443, w30444, w30445, w30446, w30447, w30448, w30449, w30450, w30451, w30452, w30453, w30454, w30455, w30456, w30457, w30458, w30459, w30460, w30461, w30462, w30463, w30464, w30465, w30466, w30467, w30468, w30469, w30470, w30471, w30472, w30473, w30474, w30475, w30476, w30477, w30478, w30479, w30480, w30481, w30482, w30483, w30484, w30485, w30486, w30487, w30488, w30489, w30490, w30491, w30492, w30493, w30494, w30495, w30496, w30497, w30498, w30499, w30500, w30501, w30502, w30503, w30504, w30505, w30506, w30507, w30508, w30509, w30510, w30511, w30512, w30513, w30514, w30515, w30516, w30517, w30518, w30519, w30520, w30521, w30522, w30523, w30524, w30525, w30526, w30527, w30528, w30529, w30530, w30531, w30532, w30533, w30534, w30535, w30536, w30537, w30538, w30539, w30540, w30541, w30542, w30543, w30544, w30545, w30546, w30547, w30548, w30549, w30550, w30551, w30552, w30553, w30554, w30555, w30556, w30557, w30558, w30559, w30560, w30561, w30562, w30563, w30564, w30565, w30566, w30567, w30568, w30569, w30570, w30571, w30572, w30573, w30574, w30575, w30576, w30577, w30578, w30579, w30580, w30581, w30582, w30583, w30584, w30585, w30586, w30587, w30588, w30589, w30590, w30591, w30592, w30593, w30594, w30595, w30596, w30597, w30598, w30599, w30600, w30601, w30602, w30603, w30604, w30605, w30606, w30607, w30608, w30609, w30610, w30611, w30612, w30613, w30614, w30615, w30616, w30617, w30618, w30619, w30620, w30621, w30622, w30623, w30624, w30625, w30626, w30627, w30628, w30629, w30630, w30631, w30632, w30633, w30634, w30635, w30636, w30637, w30638, w30639, w30640, w30641, w30642, w30643, w30644, w30645, w30646, w30647, w30648, w30649, w30650, w30651, w30652, w30653, w30654, w30655, w30656, w30657, w30658, w30659, w30660, w30661, w30662, w30663, w30664, w30665, w30666, w30667, w30668, w30669, w30670, w30671, w30672, w30673, w30674, w30675, w30676, w30677, w30678, w30679, w30680, w30681, w30682, w30683, w30684, w30685, w30686, w30687, w30688, w30689, w30690, w30691, w30692, w30693, w30694, w30695, w30696, w30697, w30698, w30699, w30700, w30701, w30702, w30703, w30704, w30705, w30706, w30707, w30708, w30709, w30710, w30711, w30712, w30713, w30714, w30715, w30716, w30717, w30718, w30719, w30720, w30721, w30722, w30723, w30724, w30725, w30726, w30727, w30728, w30729, w30730, w30731, w30732, w30733, w30734, w30735, w30736, w30737, w30738, w30739, w30740, w30741, w30742, w30743, w30744, w30745, w30746, w30747, w30748, w30749, w30750, w30751, w30752, w30753, w30754, w30755, w30756, w30757, w30758, w30759, w30760, w30761, w30762, w30763, w30764, w30765, w30766, w30767, w30768, w30769, w30770, w30771, w30772, w30773, w30774, w30775, w30776, w30777, w30778, w30779, w30780, w30781, w30782, w30783, w30784, w30785, w30786, w30787, w30788, w30789, w30790, w30791, w30792, w30793, w30794, w30795, w30796, w30797, w30798, w30799, w30800, w30801, w30802, w30803, w30804, w30805, w30806, w30807, w30808, w30809, w30810, w30811, w30812, w30813, w30814, w30815, w30816, w30817, w30818, w30819, w30820, w30821, w30822, w30823, w30824, w30825, w30826, w30827, w30828, w30829, w30830, w30831, w30832, w30833, w30834, w30835, w30836, w30837, w30838, w30839, w30840, w30841, w30842, w30843, w30844, w30845, w30846, w30847, w30848, w30849, w30850, w30851, w30852, w30853, w30854, w30855, w30856, w30857, w30858, w30859, w30860, w30861, w30862, w30863, w30864, w30865, w30866, w30867, w30868, w30869, w30870, w30871, w30872, w30873, w30874, w30875, w30876, w30877, w30878, w30879, w30880, w30881, w30882, w30883, w30884, w30885, w30886, w30887, w30888, w30889, w30890, w30891, w30892, w30893, w30894, w30895, w30896, w30897, w30898, w30899, w30900, w30901, w30902, w30903, w30904, w30905, w30906, w30907, w30908, w30909, w30910, w30911, w30912, w30913, w30914, w30915, w30916, w30917, w30918, w30919, w30920, w30921, w30922, w30923, w30924, w30925, w30926, w30927, w30928, w30929, w30930, w30931, w30932, w30933, w30934, w30935, w30936, w30937, w30938, w30939, w30940, w30941, w30942, w30943, w30944, w30945, w30946, w30947, w30948, w30949, w30950, w30951, w30952, w30953, w30954, w30955, w30956, w30957, w30958, w30959, w30960, w30961, w30962, w30963, w30964, w30965, w30966, w30967, w30968, w30969, w30970, w30971, w30972, w30973, w30974, w30975, w30976, w30977, w30978, w30979, w30980, w30981, w30982, w30983, w30984, w30985, w30986, w30987, w30988, w30989, w30990, w30991, w30992, w30993, w30994, w30995, w30996, w30997, w30998, w30999, w31000, w31001, w31002, w31003, w31004, w31005, w31006, w31007, w31008, w31009, w31010, w31011, w31012, w31013, w31014, w31015, w31016, w31017, w31018, w31019, w31020, w31021, w31022, w31023, w31024, w31025, w31026, w31027, w31028, w31029, w31030, w31031, w31032, w31033, w31034, w31035, w31036, w31037, w31038, w31039, w31040, w31041, w31042, w31043, w31044, w31045, w31046, w31047, w31048, w31049, w31050, w31051, w31052, w31053, w31054, w31055, w31056, w31057, w31058, w31059, w31060, w31061, w31062, w31063, w31064, w31065, w31066, w31067, w31068, w31069, w31070, w31071, w31072, w31073, w31074, w31075, w31076, w31077, w31078, w31079, w31080, w31081, w31082, w31083, w31084, w31085, w31086, w31087, w31088, w31089, w31090, w31091, w31092, w31093, w31094, w31095, w31096, w31097, w31098, w31099, w31100, w31101, w31102, w31103, w31104, w31105, w31106, w31107, w31108, w31109, w31110, w31111, w31112, w31113, w31114, w31115, w31116, w31117, w31118, w31119, w31120, w31121, w31122, w31123, w31124, w31125, w31126, w31127, w31128, w31129, w31130, w31131, w31132, w31133, w31134, w31135, w31136, w31137, w31138, w31139, w31140, w31141, w31142, w31143, w31144, w31145, w31146, w31147, w31148, w31149, w31150, w31151, w31152, w31153, w31154, w31155, w31156, w31157, w31158, w31159, w31160, w31161, w31162, w31163, w31164, w31165, w31166, w31167, w31168, w31169, w31170, w31171, w31172, w31173, w31174, w31175, w31176, w31177, w31178, w31179, w31180, w31181, w31182, w31183, w31184, w31185, w31186, w31187, w31188, w31189, w31190, w31191, w31192, w31193, w31194, w31195, w31196, w31197, w31198, w31199, w31200, w31201, w31202, w31203, w31204, w31205, w31206, w31207, w31208, w31209, w31210, w31211, w31212, w31213, w31214, w31215, w31216, w31217, w31218, w31219, w31220, w31221, w31222, w31223, w31224, w31225, w31226, w31227, w31228, w31229, w31230, w31231, w31232, w31233, w31234, w31235, w31236, w31237, w31238, w31239, w31240, w31241, w31242, w31243, w31244, w31245, w31246, w31247, w31248, w31249, w31250, w31251, w31252, w31253, w31254, w31255, w31256, w31257, w31258, w31259, w31260, w31261, w31262, w31263, w31264, w31265, w31266, w31267, w31268, w31269, w31270, w31271, w31272, w31273, w31274, w31275, w31276, w31277, w31278, w31279, w31280, w31281, w31282, w31283, w31284, w31285, w31286, w31287, w31288, w31289, w31290, w31291, w31292, w31293, w31294, w31295, w31296, w31297, w31298, w31299, w31300, w31301, w31302, w31303, w31304, w31305, w31306, w31307, w31308, w31309, w31310, w31311, w31312, w31313, w31314, w31315, w31316, w31317, w31318, w31319, w31320, w31321, w31322, w31323, w31324, w31325, w31326, w31327, w31328, w31329, w31330, w31331, w31332, w31333, w31334, w31335, w31336, w31337, w31338, w31339, w31340, w31341, w31342, w31343, w31344, w31345, w31346, w31347, w31348, w31349, w31350, w31351, w31352, w31353, w31354, w31355, w31356, w31357, w31358, w31359, w31360, w31361, w31362, w31363, w31364, w31365, w31366, w31367, w31368, w31369, w31370, w31371, w31372, w31373, w31374, w31375, w31376, w31377, w31378, w31379, w31380, w31381, w31382, w31383, w31384, w31385, w31386, w31387, w31388, w31389, w31390, w31391, w31392, w31393, w31394, w31395, w31396, w31397, w31398, w31399, w31400, w31401, w31402, w31403, w31404, w31405, w31406, w31407, w31408, w31409, w31410, w31411, w31412, w31413, w31414, w31415, w31416, w31417, w31418, w31419, w31420, w31421, w31422, w31423, w31424, w31425, w31426, w31427, w31428, w31429, w31430, w31431, w31432, w31433, w31434, w31435, w31436, w31437, w31438, w31439, w31440, w31441, w31442, w31443, w31444, w31445, w31446, w31447, w31448, w31449, w31450, w31451, w31452, w31453, w31454, w31455, w31456, w31457, w31458, w31459, w31460, w31461, w31462, w31463, w31464, w31465, w31466, w31467, w31468, w31469, w31470, w31471, w31472, w31473, w31474, w31475, w31476, w31477, w31478, w31479, w31480, w31481, w31482, w31483, w31484, w31485, w31486, w31487, w31488, w31489, w31490, w31491, w31492, w31493, w31494, w31495, w31496, w31497, w31498, w31499, w31500, w31501, w31502, w31503, w31504, w31505, w31506, w31507, w31508, w31509, w31510, w31511, w31512, w31513, w31514, w31515, w31516, w31517, w31518, w31519, w31520, w31521, w31522, w31523, w31524, w31525, w31526, w31527, w31528, w31529, w31530, w31531, w31532, w31533, w31534, w31535, w31536, w31537, w31538, w31539, w31540, w31541, w31542, w31543, w31544, w31545, w31546, w31547, w31548, w31549, w31550, w31551, w31552, w31553, w31554, w31555, w31556, w31557, w31558, w31559, w31560, w31561, w31562, w31563, w31564, w31565, w31566, w31567, w31568, w31569, w31570, w31571, w31572, w31573, w31574, w31575, w31576, w31577, w31578, w31579, w31580, w31581, w31582, w31583, w31584, w31585, w31586, w31587, w31588, w31589, w31590, w31591, w31592, w31593, w31594, w31595, w31596, w31597, w31598, w31599, w31600, w31601, w31602, w31603, w31604, w31605, w31606, w31607, w31608, w31609, w31610, w31611, w31612, w31613, w31614, w31615, w31616, w31617, w31618, w31619, w31620, w31621, w31622, w31623, w31624, w31625, w31626, w31627, w31628, w31629, w31630, w31631, w31632, w31633, w31634, w31635, w31636, w31637, w31638, w31639, w31640, w31641, w31642, w31643, w31644, w31645, w31646, w31647, w31648, w31649, w31650, w31651, w31652, w31653, w31654, w31655, w31656, w31657, w31658, w31659, w31660, w31661, w31662, w31663, w31664, w31665, w31666, w31667, w31668, w31669, w31670, w31671, w31672, w31673, w31674, w31675, w31676, w31677, w31678, w31679, w31680, w31681, w31682, w31683, w31684, w31685, w31686, w31687, w31688, w31689, w31690, w31691, w31692, w31693, w31694, w31695, w31696, w31697, w31698, w31699, w31700, w31701, w31702, w31703, w31704, w31705, w31706, w31707, w31708, w31709, w31710, w31711, w31712, w31713, w31714, w31715, w31716, w31717, w31718, w31719, w31720, w31721, w31722, w31723, w31724, w31725, w31726, w31727, w31728, w31729, w31730, w31731, w31732, w31733, w31734, w31735, w31736, w31737, w31738, w31739, w31740, w31741, w31742, w31743, w31744, w31745, w31746, w31747, w31748, w31749, w31750, w31751, w31752, w31753, w31754, w31755, w31756, w31757, w31758, w31759, w31760, w31761, w31762, w31763, w31764, w31765, w31766, w31767, w31768, w31769, w31770, w31771, w31772, w31773, w31774, w31775, w31776, w31777, w31778, w31779, w31780, w31781, w31782, w31783, w31784, w31785, w31786, w31787, w31788, w31789, w31790, w31791, w31792, w31793, w31794, w31795, w31796, w31797, w31798, w31799, w31800, w31801, w31802, w31803, w31804, w31805, w31806, w31807, w31808, w31809, w31810, w31811, w31812, w31813, w31814, w31815, w31816, w31817, w31818, w31819, w31820, w31821, w31822, w31823, w31824, w31825, w31826, w31827, w31828, w31829, w31830, w31831, w31832, w31833, w31834, w31835, w31836, w31837, w31838, w31839, w31840, w31841, w31842, w31843, w31844, w31845, w31846, w31847, w31848, w31849, w31850, w31851, w31852, w31853, w31854, w31855, w31856, w31857, w31858, w31859, w31860, w31861, w31862, w31863, w31864, w31865, w31866, w31867, w31868, w31869, w31870, w31871, w31872, w31873, w31874, w31875, w31876, w31877, w31878, w31879, w31880, w31881, w31882, w31883, w31884, w31885, w31886, w31887, w31888, w31889, w31890, w31891, w31892, w31893, w31894, w31895, w31896, w31897, w31898, w31899, w31900, w31901, w31902, w31903, w31904, w31905, w31906, w31907, w31908, w31909, w31910, w31911, w31912, w31913, w31914, w31915, w31916, w31917, w31918, w31919, w31920, w31921, w31922, w31923, w31924, w31925, w31926, w31927, w31928, w31929, w31930, w31931, w31932, w31933, w31934, w31935, w31936, w31937, w31938, w31939, w31940, w31941, w31942, w31943, w31944, w31945, w31946, w31947, w31948, w31949, w31950, w31951, w31952, w31953, w31954, w31955, w31956, w31957, w31958, w31959, w31960, w31961, w31962, w31963, w31964, w31965, w31966, w31967, w31968, w31969, w31970, w31971, w31972, w31973, w31974, w31975, w31976, w31977, w31978, w31979, w31980, w31981, w31982, w31983, w31984, w31985, w31986, w31987, w31988, w31989, w31990, w31991, w31992, w31993, w31994, w31995, w31996, w31997, w31998, w31999, w32000, w32001, w32002, w32003, w32004, w32005, w32006, w32007, w32008, w32009, w32010, w32011, w32012, w32013, w32014, w32015, w32016, w32017, w32018, w32019, w32020, w32021, w32022, w32023, w32024, w32025, w32026, w32027, w32028, w32029, w32030, w32031, w32032, w32033, w32034, w32035, w32036, w32037, w32038, w32039, w32040, w32041, w32042, w32043, w32044, w32045, w32046, w32047, w32048, w32049, w32050, w32051, w32052, w32053, w32054, w32055, w32056, w32057, w32058, w32059, w32060, w32061, w32062, w32063, w32064, w32065, w32066, w32067, w32068, w32069, w32070, w32071, w32072, w32073, w32074, w32075, w32076, w32077, w32078, w32079, w32080, w32081, w32082, w32083, w32084, w32085, w32086, w32087, w32088, w32089, w32090, w32091, w32092, w32093, w32094, w32095, w32096, w32097, w32098, w32099, w32100, w32101, w32102, w32103, w32104, w32105, w32106, w32107, w32108, w32109, w32110, w32111, w32112, w32113, w32114, w32115, w32116, w32117, w32118, w32119, w32120, w32121, w32122, w32123, w32124, w32125, w32126, w32127, w32128, w32129, w32130, w32131, w32132, w32133, w32134, w32135, w32136, w32137, w32138, w32139, w32140, w32141, w32142, w32143, w32144, w32145, w32146, w32147, w32148, w32149, w32150, w32151, w32152, w32153, w32154, w32155, w32156, w32157, w32158, w32159, w32160, w32161, w32162, w32163, w32164, w32165, w32166, w32167, w32168, w32169, w32170, w32171, w32172, w32173, w32174, w32175, w32176, w32177, w32178, w32179, w32180, w32181, w32182, w32183, w32184, w32185, w32186, w32187, w32188, w32189, w32190, w32191, w32192, w32193, w32194, w32195, w32196, w32197, w32198, w32199, w32200, w32201, w32202, w32203, w32204, w32205, w32206, w32207, w32208, w32209, w32210, w32211, w32212, w32213, w32214, w32215, w32216, w32217, w32218, w32219, w32220, w32221, w32222, w32223, w32224, w32225, w32226, w32227, w32228, w32229, w32230, w32231, w32232, w32233, w32234, w32235, w32236, w32237, w32238, w32239, w32240, w32241, w32242, w32243, w32244, w32245, w32246, w32247, w32248, w32249, w32250, w32251, w32252, w32253, w32254, w32255, w32256, w32257, w32258, w32259, w32260, w32261, w32262, w32263, w32264, w32265, w32266, w32267, w32268, w32269, w32270, w32271, w32272, w32273, w32274, w32275, w32276, w32277, w32278, w32279, w32280, w32281, w32282, w32283, w32284, w32285, w32286, w32287, w32288, w32289, w32290, w32291, w32292, w32293, w32294, w32295, w32296, w32297, w32298, w32299, w32300, w32301, w32302, w32303, w32304, w32305, w32306, w32307, w32308, w32309, w32310, w32311, w32312, w32313, w32314, w32315, w32316, w32317, w32318, w32319, w32320, w32321, w32322, w32323, w32324, w32325, w32326, w32327, w32328, w32329, w32330, w32331, w32332, w32333, w32334, w32335, w32336, w32337, w32338, w32339, w32340, w32341, w32342, w32343, w32344, w32345, w32346, w32347, w32348, w32349, w32350, w32351, w32352, w32353, w32354, w32355, w32356, w32357, w32358, w32359, w32360, w32361, w32362, w32363, w32364, w32365, w32366, w32367, w32368, w32369, w32370, w32371, w32372, w32373, w32374, w32375, w32376, w32377, w32378, w32379, w32380, w32381, w32382, w32383, w32384, w32385, w32386, w32387, w32388, w32389, w32390, w32391, w32392, w32393, w32394, w32395, w32396, w32397, w32398, w32399, w32400, w32401, w32402, w32403, w32404, w32405, w32406, w32407, w32408, w32409, w32410, w32411, w32412, w32413, w32414, w32415, w32416, w32417, w32418, w32419, w32420, w32421, w32422, w32423, w32424, w32425, w32426, w32427, w32428, w32429, w32430, w32431, w32432, w32433, w32434, w32435, w32436, w32437, w32438, w32439, w32440, w32441, w32442, w32443, w32444, w32445, w32446, w32447, w32448, w32449, w32450, w32451, w32452, w32453, w32454, w32455, w32456, w32457, w32458, w32459, w32460, w32461, w32462, w32463, w32464, w32465, w32466, w32467, w32468, w32469, w32470, w32471, w32472, w32473, w32474, w32475, w32476, w32477, w32478, w32479, w32480, w32481, w32482, w32483, w32484, w32485, w32486, w32487, w32488, w32489, w32490, w32491, w32492, w32493, w32494, w32495, w32496, w32497, w32498, w32499, w32500, w32501, w32502, w32503, w32504, w32505, w32506, w32507, w32508, w32509, w32510, w32511, w32512, w32513, w32514, w32515, w32516, w32517, w32518, w32519, w32520, w32521, w32522, w32523, w32524, w32525, w32526, w32527, w32528, w32529, w32530, w32531, w32532, w32533, w32534, w32535, w32536, w32537, w32538, w32539, w32540, w32541, w32542, w32543, w32544, w32545, w32546, w32547, w32548, w32549, w32550, w32551, w32552, w32553, w32554, w32555, w32556, w32557, w32558, w32559, w32560, w32561, w32562, w32563, w32564, w32565, w32566, w32567, w32568, w32569, w32570, w32571, w32572, w32573, w32574, w32575, w32576, w32577, w32578, w32579, w32580, w32581, w32582, w32583, w32584, w32585, w32586, w32587, w32588, w32589, w32590, w32591, w32592, w32593, w32594, w32595, w32596, w32597, w32598, w32599, w32600, w32601, w32602, w32603, w32604, w32605, w32606, w32607, w32608, w32609, w32610, w32611, w32612, w32613, w32614, w32615, w32616, w32617, w32618, w32619, w32620, w32621, w32622, w32623, w32624, w32625, w32626, w32627, w32628, w32629, w32630, w32631, w32632, w32633, w32634, w32635, w32636, w32637, w32638, w32639, w32640, w32641, w32642, w32643, w32644, w32645, w32646, w32647, w32648, w32649, w32650, w32651, w32652, w32653, w32654, w32655, w32656, w32657, w32658, w32659, w32660, w32661, w32662, w32663, w32664, w32665, w32666, w32667, w32668, w32669, w32670, w32671, w32672, w32673, w32674, w32675, w32676, w32677, w32678, w32679, w32680, w32681, w32682, w32683, w32684, w32685, w32686, w32687, w32688, w32689, w32690, w32691, w32692, w32693, w32694, w32695, w32696, w32697, w32698, w32699, w32700, w32701, w32702, w32703, w32704, w32705, w32706, w32707, w32708, w32709, w32710, w32711, w32712, w32713, w32714, w32715, w32716, w32717, w32718, w32719, w32720, w32721, w32722, w32723, w32724, w32725, w32726, w32727, w32728, w32729, w32730, w32731, w32732, w32733, w32734, w32735, w32736, w32737, w32738, w32739, w32740, w32741, w32742, w32743, w32744, w32745, w32746, w32747, w32748, w32749, w32750, w32751, w32752, w32753, w32754, w32755, w32756, w32757, w32758, w32759, w32760, w32761, w32762, w32763, w32764, w32765, w32766, w32767, w32768, w32769, w32770, w32771, w32772, w32773, w32774, w32775, w32776, w32777, w32778, w32779, w32780, w32781, w32782, w32783, w32784, w32785, w32786, w32787, w32788, w32789, w32790, w32791, w32792, w32793, w32794, w32795, w32796, w32797, w32798, w32799, w32800, w32801, w32802, w32803, w32804, w32805, w32806, w32807, w32808, w32809, w32810, w32811, w32812, w32813, w32814, w32815, w32816, w32817, w32818, w32819, w32820, w32821, w32822, w32823, w32824, w32825, w32826, w32827, w32828, w32829, w32830, w32831, w32832, w32833, w32834, w32835, w32836, w32837, w32838, w32839, w32840, w32841, w32842, w32843, w32844, w32845, w32846, w32847, w32848, w32849, w32850, w32851, w32852, w32853, w32854, w32855, w32856, w32857, w32858, w32859, w32860, w32861, w32862, w32863, w32864, w32865, w32866, w32867, w32868, w32869, w32870, w32871, w32872, w32873, w32874, w32875, w32876, w32877, w32878, w32879, w32880, w32881, w32882, w32883, w32884, w32885, w32886, w32887, w32888, w32889, w32890, w32891, w32892, w32893, w32894, w32895, w32896, w32897, w32898, w32899, w32900, w32901, w32902, w32903, w32904, w32905, w32906, w32907, w32908, w32909, w32910, w32911, w32912, w32913, w32914, w32915, w32916, w32917, w32918, w32919, w32920, w32921, w32922, w32923, w32924, w32925, w32926, w32927, w32928, w32929, w32930, w32931, w32932, w32933, w32934, w32935, w32936, w32937, w32938, w32939, w32940, w32941, w32942, w32943, w32944, w32945, w32946, w32947, w32948, w32949, w32950, w32951, w32952, w32953, w32954, w32955, w32956, w32957, w32958, w32959, w32960, w32961, w32962, w32963, w32964, w32965, w32966, w32967, w32968, w32969, w32970, w32971, w32972, w32973, w32974, w32975, w32976, w32977, w32978, w32979, w32980, w32981, w32982, w32983, w32984, w32985, w32986, w32987, w32988, w32989, w32990, w32991, w32992, w32993, w32994, w32995, w32996, w32997, w32998, w32999, w33000, w33001, w33002, w33003, w33004, w33005, w33006, w33007, w33008, w33009, w33010, w33011, w33012, w33013, w33014, w33015, w33016, w33017, w33018, w33019, w33020, w33021, w33022, w33023, w33024, w33025, w33026, w33027, w33028, w33029, w33030, w33031, w33032, w33033, w33034, w33035, w33036, w33037, w33038, w33039, w33040, w33041, w33042, w33043, w33044, w33045, w33046, w33047, w33048, w33049, w33050, w33051, w33052, w33053, w33054, w33055, w33056, w33057, w33058, w33059, w33060, w33061, w33062, w33063, w33064, w33065, w33066, w33067, w33068, w33069, w33070, w33071, w33072, w33073, w33074, w33075, w33076, w33077, w33078, w33079, w33080, w33081, w33082, w33083, w33084, w33085, w33086, w33087, w33088, w33089, w33090, w33091, w33092, w33093, w33094, w33095, w33096, w33097, w33098, w33099, w33100, w33101, w33102, w33103, w33104, w33105, w33106, w33107, w33108, w33109, w33110, w33111, w33112, w33113, w33114, w33115, w33116, w33117, w33118, w33119, w33120, w33121, w33122, w33123, w33124, w33125, w33126, w33127, w33128, w33129, w33130, w33131, w33132, w33133, w33134, w33135, w33136, w33137, w33138, w33139, w33140, w33141, w33142, w33143, w33144, w33145, w33146, w33147, w33148, w33149, w33150, w33151, w33152, w33153, w33154, w33155, w33156, w33157, w33158, w33159, w33160, w33161, w33162, w33163, w33164, w33165, w33166, w33167, w33168, w33169, w33170, w33171, w33172, w33173, w33174, w33175, w33176, w33177, w33178, w33179, w33180, w33181, w33182, w33183, w33184, w33185, w33186, w33187, w33188, w33189, w33190, w33191, w33192, w33193, w33194, w33195, w33196, w33197, w33198, w33199, w33200, w33201, w33202, w33203, w33204, w33205, w33206, w33207, w33208, w33209, w33210, w33211, w33212, w33213, w33214, w33215, w33216, w33217, w33218, w33219, w33220, w33221, w33222, w33223, w33224, w33225, w33226, w33227, w33228, w33229, w33230, w33231, w33232, w33233, w33234, w33235, w33236, w33237, w33238, w33239, w33240, w33241, w33242, w33243, w33244, w33245, w33246, w33247, w33248, w33249, w33250, w33251, w33252, w33253, w33254, w33255, w33256, w33257, w33258, w33259, w33260, w33261, w33262, w33263, w33264, w33265, w33266, w33267, w33268, w33269, w33270, w33271, w33272, w33273, w33274, w33275, w33276, w33277, w33278, w33279, w33280, w33281, w33282, w33283, w33284, w33285, w33286, w33287, w33288, w33289, w33290, w33291, w33292, w33293, w33294, w33295, w33296, w33297, w33298, w33299, w33300, w33301, w33302, w33303, w33304, w33305, w33306, w33307, w33308, w33309, w33310, w33311, w33312, w33313, w33314, w33315, w33316, w33317, w33318, w33319, w33320, w33321, w33322, w33323, w33324, w33325, w33326, w33327, w33328, w33329, w33330, w33331, w33332, w33333, w33334, w33335, w33336, w33337, w33338, w33339, w33340, w33341, w33342, w33343, w33344, w33345, w33346, w33347, w33348, w33349, w33350, w33351, w33352, w33353, w33354, w33355, w33356, w33357, w33358, w33359, w33360, w33361, w33362, w33363, w33364, w33365, w33366, w33367, w33368, w33369, w33370, w33371, w33372, w33373, w33374, w33375, w33376, w33377, w33378, w33379, w33380, w33381, w33382, w33383, w33384, w33385, w33386, w33387, w33388, w33389, w33390, w33391, w33392, w33393, w33394, w33395, w33396, w33397, w33398, w33399, w33400, w33401, w33402, w33403, w33404, w33405, w33406, w33407, w33408, w33409, w33410, w33411, w33412, w33413, w33414, w33415, w33416, w33417, w33418, w33419, w33420, w33421, w33422, w33423, w33424, w33425, w33426, w33427, w33428, w33429, w33430, w33431, w33432, w33433, w33434, w33435, w33436, w33437, w33438, w33439, w33440, w33441, w33442, w33443, w33444, w33445, w33446, w33447, w33448, w33449, w33450, w33451, w33452, w33453, w33454, w33455, w33456, w33457, w33458, w33459, w33460, w33461, w33462, w33463, w33464, w33465, w33466, w33467, w33468, w33469, w33470, w33471, w33472, w33473, w33474, w33475, w33476, w33477, w33478, w33479, w33480, w33481, w33482, w33483, w33484, w33485, w33486, w33487, w33488, w33489, w33490, w33491, w33492, w33493, w33494, w33495, w33496, w33497, w33498, w33499, w33500, w33501, w33502, w33503, w33504, w33505, w33506, w33507, w33508, w33509, w33510, w33511, w33512, w33513, w33514, w33515, w33516, w33517, w33518, w33519, w33520, w33521, w33522, w33523, w33524, w33525, w33526, w33527, w33528, w33529, w33530, w33531, w33532, w33533, w33534, w33535, w33536, w33537, w33538, w33539, w33540, w33541, w33542, w33543, w33544, w33545, w33546, w33547, w33548, w33549, w33550, w33551, w33552, w33553, w33554, w33555, w33556, w33557, w33558, w33559, w33560, w33561, w33562, w33563, w33564, w33565, w33566, w33567, w33568, w33569, w33570, w33571, w33572, w33573, w33574, w33575, w33576, w33577, w33578, w33579, w33580, w33581, w33582, w33583, w33584, w33585, w33586, w33587, w33588, w33589, w33590, w33591, w33592, w33593, w33594, w33595, w33596, w33597, w33598, w33599, w33600, w33601, w33602, w33603, w33604, w33605, w33606, w33607, w33608, w33609, w33610, w33611, w33612, w33613, w33614, w33615, w33616, w33617, w33618, w33619, w33620, w33621, w33622, w33623, w33624, w33625, w33626, w33627, w33628, w33629, w33630, w33631, w33632, w33633, w33634, w33635, w33636, w33637, w33638, w33639, w33640, w33641, w33642, w33643, w33644, w33645, w33646, w33647, w33648, w33649, w33650, w33651, w33652, w33653, w33654, w33655, w33656, w33657, w33658, w33659, w33660, w33661, w33662, w33663, w33664, w33665, w33666, w33667, w33668, w33669, w33670, w33671, w33672, w33673, w33674, w33675, w33676, w33677, w33678, w33679, w33680, w33681, w33682, w33683, w33684, w33685, w33686, w33687, w33688, w33689, w33690, w33691, w33692, w33693, w33694, w33695, w33696, w33697, w33698, w33699, w33700, w33701, w33702, w33703, w33704, w33705, w33706, w33707, w33708, w33709, w33710, w33711, w33712, w33713, w33714, w33715, w33716, w33717, w33718, w33719, w33720, w33721, w33722, w33723, w33724, w33725, w33726, w33727, w33728, w33729, w33730, w33731, w33732, w33733, w33734, w33735, w33736, w33737, w33738, w33739, w33740, w33741, w33742, w33743, w33744, w33745, w33746, w33747, w33748, w33749, w33750, w33751, w33752, w33753, w33754, w33755, w33756, w33757, w33758, w33759, w33760, w33761, w33762, w33763, w33764, w33765, w33766, w33767, w33768, w33769, w33770, w33771, w33772, w33773, w33774, w33775, w33776, w33777, w33778, w33779, w33780, w33781, w33782, w33783, w33784, w33785, w33786, w33787, w33788, w33789, w33790, w33791, w33792, w33793, w33794, w33795, w33796, w33797, w33798, w33799, w33800, w33801, w33802, w33803, w33804, w33805, w33806, w33807, w33808, w33809, w33810, w33811, w33812, w33813, w33814, w33815, w33816, w33817, w33818, w33819, w33820, w33821, w33822, w33823, w33824, w33825, w33826, w33827, w33828, w33829, w33830, w33831, w33832, w33833, w33834, w33835, w33836, w33837, w33838, w33839, w33840, w33841, w33842, w33843, w33844, w33845, w33846, w33847, w33848, w33849, w33850, w33851, w33852, w33853, w33854, w33855, w33856, w33857, w33858, w33859, w33860, w33861, w33862, w33863, w33864, w33865, w33866, w33867, w33868, w33869, w33870, w33871, w33872, w33873, w33874, w33875, w33876, w33877, w33878, w33879, w33880, w33881, w33882, w33883, w33884, w33885, w33886, w33887, w33888, w33889, w33890, w33891, w33892, w33893, w33894, w33895, w33896, w33897, w33898, w33899, w33900, w33901, w33902, w33903, w33904, w33905, w33906, w33907, w33908, w33909, w33910, w33911, w33912, w33913, w33914, w33915, w33916, w33917, w33918, w33919, w33920, w33921, w33922, w33923, w33924, w33925, w33926, w33927, w33928, w33929, w33930, w33931, w33932, w33933, w33934, w33935, w33936, w33937, w33938, w33939, w33940, w33941, w33942, w33943, w33944, w33945, w33946, w33947, w33948, w33949, w33950, w33951, w33952, w33953, w33954, w33955, w33956, w33957, w33958, w33959, w33960, w33961, w33962, w33963, w33964, w33965, w33966, w33967, w33968, w33969, w33970, w33971, w33972, w33973, w33974, w33975, w33976, w33977, w33978, w33979, w33980, w33981, w33982, w33983, w33984, w33985, w33986, w33987, w33988, w33989, w33990, w33991, w33992, w33993, w33994, w33995, w33996, w33997, w33998, w33999, w34000, w34001, w34002, w34003, w34004, w34005, w34006, w34007, w34008, w34009, w34010, w34011, w34012, w34013, w34014, w34015, w34016, w34017, w34018, w34019, w34020, w34021, w34022, w34023, w34024, w34025, w34026, w34027, w34028, w34029, w34030, w34031, w34032, w34033, w34034, w34035, w34036, w34037, w34038, w34039, w34040, w34041, w34042, w34043, w34044, w34045, w34046, w34047, w34048, w34049, w34050, w34051, w34052, w34053, w34054, w34055, w34056, w34057, w34058, w34059, w34060, w34061, w34062, w34063, w34064, w34065, w34066, w34067, w34068, w34069, w34070, w34071, w34072, w34073, w34074, w34075, w34076, w34077, w34078, w34079, w34080, w34081, w34082, w34083, w34084, w34085, w34086, w34087, w34088, w34089, w34090, w34091, w34092, w34093, w34094, w34095, w34096, w34097, w34098, w34099, w34100, w34101, w34102, w34103, w34104, w34105, w34106, w34107, w34108, w34109, w34110, w34111, w34112, w34113, w34114, w34115, w34116, w34117, w34118, w34119, w34120, w34121, w34122, w34123, w34124, w34125, w34126, w34127, w34128, w34129, w34130, w34131, w34132, w34133, w34134, w34135, w34136, w34137, w34138, w34139, w34140, w34141, w34142, w34143, w34144, w34145, w34146, w34147, w34148, w34149, w34150, w34151, w34152, w34153, w34154, w34155, w34156, w34157, w34158, w34159, w34160, w34161, w34162, w34163, w34164, w34165, w34166, w34167, w34168, w34169, w34170, w34171, w34172, w34173, w34174, w34175, w34176, w34177, w34178, w34179, w34180, w34181, w34182, w34183, w34184, w34185, w34186, w34187, w34188, w34189, w34190, w34191, w34192, w34193, w34194, w34195, w34196, w34197, w34198, w34199, w34200, w34201, w34202, w34203, w34204, w34205, w34206, w34207, w34208, w34209, w34210, w34211, w34212, w34213, w34214, w34215, w34216, w34217, w34218, w34219, w34220, w34221, w34222, w34223, w34224, w34225, w34226, w34227, w34228, w34229, w34230, w34231, w34232, w34233, w34234, w34235, w34236, w34237, w34238, w34239, w34240, w34241, w34242, w34243, w34244, w34245, w34246, w34247, w34248, w34249, w34250, w34251, w34252, w34253, w34254, w34255, w34256, w34257, w34258, w34259, w34260, w34261, w34262, w34263, w34264, w34265, w34266, w34267, w34268, w34269, w34270, w34271, w34272, w34273, w34274, w34275, w34276, w34277, w34278, w34279, w34280, w34281, w34282, w34283, w34284, w34285, w34286, w34287, w34288, w34289, w34290, w34291, w34292, w34293, w34294, w34295, w34296, w34297, w34298, w34299, w34300, w34301, w34302, w34303, w34304, w34305, w34306, w34307, w34308, w34309, w34310, w34311, w34312, w34313, w34314, w34315, w34316, w34317, w34318, w34319, w34320, w34321, w34322, w34323, w34324, w34325, w34326, w34327, w34328, w34329, w34330, w34331, w34332, w34333, w34334, w34335, w34336, w34337, w34338, w34339, w34340, w34341, w34342, w34343, w34344, w34345, w34346, w34347, w34348, w34349, w34350, w34351, w34352, w34353, w34354, w34355, w34356, w34357, w34358, w34359, w34360, w34361, w34362, w34363, w34364, w34365, w34366, w34367, w34368, w34369, w34370, w34371, w34372, w34373, w34374, w34375, w34376, w34377, w34378, w34379, w34380, w34381, w34382, w34383, w34384, w34385, w34386, w34387, w34388, w34389, w34390, w34391, w34392, w34393, w34394, w34395, w34396, w34397, w34398, w34399, w34400, w34401, w34402, w34403, w34404, w34405, w34406, w34407, w34408, w34409, w34410, w34411, w34412, w34413, w34414, w34415, w34416, w34417, w34418, w34419, w34420, w34421, w34422, w34423, w34424, w34425, w34426, w34427, w34428, w34429, w34430, w34431, w34432, w34433, w34434, w34435, w34436, w34437, w34438, w34439, w34440, w34441, w34442, w34443, w34444, w34445, w34446, w34447, w34448, w34449, w34450, w34451, w34452, w34453, w34454, w34455, w34456, w34457, w34458, w34459, w34460, w34461, w34462, w34463, w34464, w34465, w34466, w34467, w34468, w34469, w34470, w34471, w34472, w34473, w34474, w34475, w34476, w34477, w34478, w34479, w34480, w34481, w34482, w34483, w34484, w34485, w34486, w34487, w34488, w34489, w34490, w34491, w34492, w34493, w34494, w34495, w34496, w34497, w34498, w34499, w34500, w34501, w34502, w34503, w34504, w34505, w34506, w34507, w34508, w34509, w34510, w34511, w34512, w34513, w34514, w34515, w34516, w34517, w34518, w34519, w34520, w34521, w34522, w34523, w34524, w34525, w34526, w34527, w34528, w34529, w34530, w34531, w34532, w34533, w34534, w34535, w34536, w34537, w34538, w34539, w34540, w34541, w34542, w34543, w34544, w34545, w34546, w34547, w34548, w34549, w34550, w34551, w34552, w34553, w34554, w34555, w34556, w34557, w34558, w34559, w34560, w34561, w34562, w34563, w34564, w34565, w34566, w34567, w34568, w34569, w34570, w34571, w34572, w34573, w34574, w34575, w34576, w34577, w34578, w34579, w34580, w34581, w34582, w34583, w34584, w34585, w34586, w34587, w34588, w34589, w34590, w34591, w34592, w34593, w34594, w34595, w34596, w34597, w34598, w34599, w34600, w34601, w34602, w34603, w34604, w34605, w34606, w34607, w34608, w34609, w34610, w34611, w34612, w34613, w34614, w34615, w34616, w34617, w34618, w34619, w34620, w34621, w34622, w34623, w34624, w34625, w34626, w34627, w34628, w34629, w34630, w34631, w34632, w34633, w34634, w34635, w34636, w34637, w34638, w34639, w34640, w34641, w34642, w34643, w34644, w34645, w34646, w34647, w34648, w34649, w34650, w34651, w34652, w34653, w34654, w34655, w34656, w34657, w34658, w34659, w34660, w34661, w34662, w34663, w34664, w34665, w34666, w34667, w34668, w34669, w34670, w34671, w34672, w34673, w34674, w34675, w34676, w34677, w34678, w34679, w34680, w34681, w34682, w34683, w34684, w34685, w34686, w34687, w34688, w34689, w34690, w34691, w34692, w34693, w34694, w34695, w34696, w34697, w34698, w34699, w34700, w34701, w34702, w34703, w34704, w34705, w34706, w34707, w34708, w34709, w34710, w34711, w34712, w34713, w34714, w34715, w34716, w34717, w34718, w34719, w34720, w34721, w34722, w34723, w34724, w34725, w34726, w34727, w34728, w34729, w34730, w34731, w34732, w34733, w34734, w34735, w34736, w34737, w34738, w34739, w34740, w34741, w34742, w34743, w34744, w34745, w34746, w34747, w34748, w34749, w34750, w34751, w34752, w34753, w34754, w34755, w34756, w34757, w34758, w34759, w34760, w34761, w34762, w34763, w34764, w34765, w34766, w34767, w34768, w34769, w34770, w34771, w34772, w34773, w34774, w34775, w34776, w34777, w34778, w34779, w34780, w34781, w34782, w34783, w34784, w34785, w34786, w34787, w34788, w34789, w34790, w34791, w34792, w34793, w34794, w34795, w34796, w34797, w34798, w34799, w34800, w34801, w34802, w34803, w34804, w34805, w34806, w34807, w34808, w34809, w34810, w34811, w34812, w34813, w34814, w34815, w34816, w34817, w34818, w34819, w34820, w34821, w34822, w34823, w34824, w34825, w34826, w34827, w34828, w34829, w34830, w34831, w34832, w34833, w34834, w34835, w34836, w34837, w34838, w34839, w34840, w34841, w34842, w34843, w34844, w34845, w34846, w34847, w34848, w34849, w34850, w34851, w34852, w34853, w34854, w34855, w34856, w34857, w34858, w34859, w34860, w34861, w34862, w34863, w34864, w34865, w34866, w34867, w34868, w34869, w34870, w34871, w34872, w34873, w34874, w34875, w34876, w34877, w34878, w34879, w34880, w34881, w34882, w34883, w34884, w34885, w34886, w34887, w34888, w34889, w34890, w34891, w34892, w34893, w34894, w34895, w34896, w34897, w34898, w34899, w34900, w34901, w34902, w34903, w34904, w34905, w34906, w34907, w34908, w34909, w34910, w34911, w34912, w34913, w34914, w34915, w34916, w34917, w34918, w34919, w34920, w34921, w34922, w34923, w34924, w34925, w34926, w34927, w34928, w34929, w34930, w34931, w34932, w34933, w34934, w34935, w34936, w34937, w34938, w34939, w34940, w34941, w34942, w34943, w34944, w34945, w34946, w34947, w34948, w34949, w34950, w34951, w34952, w34953, w34954, w34955, w34956, w34957, w34958, w34959, w34960, w34961, w34962, w34963, w34964, w34965, w34966, w34967, w34968, w34969, w34970, w34971, w34972, w34973, w34974, w34975, w34976, w34977, w34978, w34979, w34980, w34981, w34982, w34983, w34984, w34985, w34986, w34987, w34988, w34989, w34990, w34991, w34992, w34993, w34994, w34995, w34996, w34997, w34998, w34999, w35000, w35001, w35002, w35003, w35004, w35005, w35006, w35007, w35008, w35009, w35010, w35011, w35012, w35013, w35014, w35015, w35016, w35017, w35018, w35019, w35020, w35021, w35022, w35023, w35024, w35025, w35026, w35027, w35028, w35029, w35030, w35031, w35032, w35033, w35034, w35035, w35036, w35037, w35038, w35039, w35040, w35041, w35042, w35043, w35044, w35045, w35046, w35047, w35048, w35049, w35050, w35051, w35052, w35053, w35054, w35055, w35056, w35057, w35058, w35059, w35060, w35061, w35062, w35063, w35064, w35065, w35066, w35067, w35068, w35069, w35070, w35071, w35072, w35073, w35074, w35075, w35076, w35077, w35078, w35079, w35080, w35081, w35082, w35083, w35084, w35085, w35086, w35087, w35088, w35089, w35090, w35091, w35092, w35093, w35094, w35095, w35096, w35097, w35098, w35099, w35100, w35101, w35102, w35103, w35104, w35105, w35106, w35107, w35108, w35109, w35110, w35111, w35112, w35113, w35114, w35115, w35116, w35117, w35118, w35119, w35120, w35121, w35122, w35123, w35124, w35125, w35126, w35127, w35128, w35129, w35130, w35131, w35132, w35133, w35134, w35135, w35136, w35137, w35138, w35139, w35140, w35141, w35142, w35143, w35144, w35145, w35146, w35147, w35148, w35149, w35150, w35151, w35152, w35153, w35154, w35155, w35156, w35157, w35158, w35159, w35160, w35161, w35162, w35163, w35164, w35165, w35166, w35167, w35168, w35169, w35170, w35171, w35172, w35173, w35174, w35175, w35176, w35177, w35178, w35179, w35180, w35181, w35182, w35183, w35184, w35185, w35186, w35187, w35188, w35189, w35190, w35191, w35192, w35193, w35194, w35195, w35196, w35197, w35198, w35199, w35200, w35201, w35202, w35203, w35204, w35205, w35206, w35207, w35208, w35209, w35210, w35211, w35212, w35213, w35214, w35215, w35216, w35217, w35218, w35219, w35220, w35221, w35222, w35223, w35224, w35225, w35226, w35227, w35228, w35229, w35230, w35231, w35232, w35233, w35234, w35235, w35236, w35237, w35238, w35239, w35240, w35241, w35242, w35243, w35244, w35245, w35246, w35247, w35248, w35249, w35250, w35251, w35252, w35253, w35254, w35255, w35256, w35257, w35258, w35259, w35260, w35261, w35262, w35263, w35264, w35265, w35266, w35267, w35268, w35269, w35270, w35271, w35272, w35273, w35274, w35275, w35276, w35277, w35278, w35279, w35280, w35281, w35282, w35283, w35284, w35285, w35286, w35287, w35288, w35289, w35290, w35291, w35292, w35293, w35294, w35295, w35296, w35297, w35298, w35299, w35300, w35301, w35302, w35303, w35304, w35305, w35306, w35307, w35308, w35309, w35310, w35311, w35312, w35313, w35314, w35315, w35316, w35317, w35318, w35319, w35320, w35321, w35322, w35323, w35324, w35325, w35326, w35327, w35328, w35329, w35330, w35331, w35332, w35333, w35334, w35335, w35336, w35337, w35338, w35339, w35340, w35341, w35342, w35343, w35344, w35345, w35346, w35347, w35348, w35349, w35350, w35351, w35352, w35353, w35354, w35355, w35356, w35357, w35358, w35359, w35360, w35361, w35362, w35363, w35364, w35365, w35366, w35367, w35368, w35369, w35370, w35371, w35372, w35373, w35374, w35375, w35376, w35377, w35378, w35379, w35380, w35381, w35382, w35383, w35384, w35385, w35386, w35387, w35388, w35389, w35390, w35391, w35392, w35393, w35394, w35395, w35396, w35397, w35398, w35399, w35400, w35401, w35402, w35403, w35404, w35405, w35406, w35407, w35408, w35409, w35410, w35411, w35412, w35413, w35414, w35415, w35416, w35417, w35418, w35419, w35420, w35421, w35422, w35423, w35424, w35425, w35426, w35427, w35428, w35429, w35430, w35431, w35432, w35433, w35434, w35435, w35436, w35437, w35438, w35439, w35440, w35441, w35442, w35443, w35444, w35445, w35446, w35447, w35448, w35449, w35450, w35451, w35452, w35453, w35454, w35455, w35456, w35457, w35458, w35459, w35460, w35461, w35462, w35463, w35464, w35465, w35466, w35467, w35468, w35469, w35470, w35471, w35472, w35473, w35474, w35475, w35476, w35477, w35478, w35479, w35480, w35481, w35482, w35483, w35484, w35485, w35486, w35487, w35488, w35489, w35490, w35491, w35492, w35493, w35494, w35495, w35496, w35497, w35498, w35499, w35500, w35501, w35502, w35503, w35504, w35505, w35506, w35507, w35508, w35509, w35510, w35511, w35512, w35513, w35514, w35515, w35516, w35517, w35518, w35519, w35520, w35521, w35522, w35523, w35524, w35525, w35526, w35527, w35528, w35529, w35530, w35531, w35532, w35533, w35534, w35535, w35536, w35537, w35538, w35539, w35540, w35541, w35542, w35543, w35544, w35545, w35546, w35547, w35548, w35549, w35550, w35551, w35552, w35553, w35554, w35555, w35556, w35557, w35558, w35559, w35560, w35561, w35562, w35563, w35564, w35565, w35566, w35567, w35568, w35569, w35570, w35571, w35572, w35573, w35574, w35575, w35576, w35577, w35578, w35579, w35580, w35581, w35582, w35583, w35584, w35585, w35586, w35587, w35588, w35589, w35590, w35591, w35592, w35593, w35594, w35595, w35596, w35597, w35598, w35599, w35600, w35601, w35602, w35603, w35604, w35605, w35606, w35607, w35608, w35609, w35610, w35611, w35612, w35613, w35614, w35615, w35616, w35617, w35618, w35619, w35620, w35621, w35622, w35623, w35624, w35625, w35626, w35627, w35628, w35629, w35630, w35631, w35632, w35633, w35634, w35635, w35636, w35637, w35638, w35639, w35640, w35641, w35642, w35643, w35644, w35645, w35646, w35647, w35648, w35649, w35650, w35651, w35652, w35653, w35654, w35655, w35656, w35657, w35658, w35659, w35660, w35661, w35662, w35663, w35664, w35665, w35666, w35667, w35668, w35669, w35670, w35671, w35672, w35673, w35674, w35675, w35676, w35677, w35678, w35679, w35680, w35681, w35682, w35683, w35684, w35685, w35686, w35687, w35688, w35689, w35690, w35691, w35692, w35693, w35694, w35695, w35696, w35697, w35698, w35699, w35700, w35701, w35702, w35703, w35704, w35705, w35706, w35707, w35708, w35709, w35710, w35711, w35712, w35713, w35714, w35715, w35716, w35717, w35718, w35719, w35720, w35721, w35722, w35723, w35724, w35725, w35726, w35727, w35728, w35729, w35730, w35731, w35732, w35733, w35734, w35735, w35736, w35737, w35738, w35739, w35740, w35741, w35742, w35743, w35744, w35745, w35746, w35747, w35748, w35749, w35750, w35751, w35752, w35753, w35754, w35755, w35756, w35757, w35758, w35759, w35760, w35761, w35762, w35763, w35764, w35765, w35766, w35767, w35768, w35769, w35770, w35771, w35772, w35773, w35774, w35775, w35776, w35777, w35778, w35779, w35780, w35781, w35782, w35783, w35784, w35785, w35786, w35787, w35788, w35789, w35790, w35791, w35792, w35793, w35794, w35795, w35796, w35797, w35798, w35799, w35800, w35801, w35802, w35803, w35804, w35805, w35806, w35807, w35808, w35809, w35810, w35811, w35812, w35813, w35814, w35815, w35816, w35817, w35818, w35819, w35820, w35821, w35822, w35823, w35824, w35825, w35826, w35827, w35828, w35829, w35830, w35831, w35832, w35833, w35834, w35835, w35836, w35837, w35838, w35839, w35840, w35841, w35842, w35843, w35844, w35845, w35846, w35847, w35848, w35849, w35850, w35851, w35852, w35853, w35854, w35855, w35856, w35857, w35858, w35859, w35860, w35861, w35862, w35863, w35864, w35865, w35866, w35867, w35868, w35869, w35870, w35871, w35872, w35873, w35874, w35875, w35876, w35877, w35878, w35879, w35880, w35881, w35882, w35883, w35884, w35885, w35886, w35887, w35888, w35889, w35890, w35891, w35892, w35893, w35894, w35895, w35896, w35897, w35898, w35899, w35900, w35901, w35902, w35903, w35904, w35905, w35906, w35907, w35908, w35909, w35910, w35911, w35912, w35913, w35914, w35915, w35916, w35917, w35918, w35919, w35920, w35921, w35922, w35923, w35924, w35925, w35926, w35927, w35928, w35929, w35930, w35931, w35932, w35933, w35934, w35935, w35936, w35937, w35938, w35939, w35940, w35941, w35942, w35943, w35944, w35945, w35946, w35947, w35948, w35949, w35950, w35951, w35952, w35953, w35954, w35955, w35956, w35957, w35958, w35959, w35960, w35961, w35962, w35963, w35964, w35965, w35966, w35967, w35968, w35969, w35970, w35971, w35972, w35973, w35974, w35975, w35976, w35977, w35978, w35979, w35980, w35981, w35982, w35983, w35984, w35985, w35986, w35987, w35988, w35989, w35990, w35991, w35992, w35993, w35994, w35995, w35996, w35997, w35998, w35999, w36000, w36001, w36002, w36003, w36004, w36005, w36006, w36007, w36008, w36009, w36010, w36011, w36012, w36013, w36014, w36015, w36016, w36017, w36018, w36019, w36020, w36021, w36022, w36023, w36024, w36025, w36026, w36027, w36028, w36029, w36030, w36031, w36032, w36033, w36034, w36035, w36036, w36037, w36038, w36039, w36040, w36041, w36042, w36043, w36044, w36045, w36046, w36047, w36048, w36049, w36050, w36051, w36052, w36053, w36054, w36055, w36056, w36057, w36058, w36059, w36060, w36061, w36062, w36063, w36064, w36065, w36066, w36067, w36068, w36069, w36070, w36071, w36072, w36073, w36074, w36075, w36076, w36077, w36078, w36079, w36080, w36081, w36082, w36083, w36084, w36085, w36086, w36087, w36088, w36089, w36090, w36091, w36092, w36093, w36094, w36095, w36096, w36097, w36098, w36099, w36100, w36101, w36102, w36103, w36104, w36105, w36106, w36107, w36108, w36109, w36110, w36111, w36112, w36113, w36114, w36115, w36116, w36117, w36118, w36119, w36120, w36121, w36122, w36123, w36124, w36125, w36126, w36127, w36128, w36129, w36130, w36131, w36132, w36133, w36134, w36135, w36136, w36137, w36138, w36139, w36140, w36141, w36142, w36143, w36144, w36145, w36146, w36147, w36148, w36149, w36150, w36151, w36152, w36153, w36154, w36155, w36156, w36157, w36158, w36159, w36160, w36161, w36162, w36163, w36164, w36165, w36166, w36167, w36168, w36169, w36170, w36171, w36172, w36173, w36174, w36175, w36176, w36177, w36178, w36179, w36180, w36181, w36182, w36183, w36184, w36185, w36186, w36187, w36188, w36189, w36190, w36191, w36192, w36193, w36194, w36195, w36196, w36197, w36198, w36199, w36200, w36201, w36202, w36203, w36204, w36205, w36206, w36207, w36208, w36209, w36210, w36211, w36212, w36213, w36214, w36215, w36216, w36217, w36218, w36219, w36220, w36221, w36222, w36223, w36224, w36225, w36226, w36227, w36228, w36229, w36230, w36231, w36232, w36233, w36234, w36235, w36236, w36237, w36238, w36239, w36240, w36241, w36242, w36243, w36244, w36245, w36246, w36247, w36248, w36249, w36250, w36251, w36252, w36253, w36254, w36255, w36256, w36257, w36258, w36259, w36260, w36261, w36262, w36263, w36264, w36265, w36266, w36267, w36268, w36269, w36270, w36271, w36272, w36273, w36274, w36275, w36276, w36277, w36278, w36279, w36280, w36281, w36282, w36283, w36284, w36285, w36286, w36287, w36288, w36289, w36290, w36291, w36292, w36293, w36294, w36295, w36296, w36297, w36298, w36299, w36300, w36301, w36302, w36303, w36304, w36305, w36306, w36307, w36308, w36309, w36310, w36311, w36312, w36313, w36314, w36315, w36316, w36317, w36318, w36319, w36320, w36321, w36322, w36323, w36324, w36325, w36326, w36327, w36328, w36329, w36330, w36331, w36332, w36333, w36334, w36335, w36336, w36337, w36338, w36339, w36340, w36341, w36342, w36343, w36344, w36345, w36346, w36347, w36348, w36349, w36350, w36351, w36352, w36353, w36354, w36355, w36356, w36357, w36358, w36359, w36360, w36361, w36362, w36363, w36364, w36365, w36366, w36367, w36368, w36369, w36370, w36371, w36372, w36373, w36374, w36375, w36376, w36377, w36378, w36379, w36380, w36381, w36382, w36383, w36384, w36385, w36386, w36387, w36388, w36389, w36390, w36391, w36392, w36393, w36394, w36395, w36396, w36397, w36398, w36399, w36400, w36401, w36402, w36403, w36404, w36405, w36406, w36407, w36408, w36409, w36410, w36411, w36412, w36413, w36414, w36415, w36416, w36417, w36418, w36419, w36420, w36421, w36422, w36423, w36424, w36425, w36426, w36427, w36428, w36429, w36430, w36431, w36432, w36433, w36434, w36435, w36436, w36437, w36438, w36439, w36440, w36441, w36442, w36443, w36444, w36445, w36446, w36447, w36448, w36449, w36450, w36451, w36452, w36453, w36454, w36455, w36456, w36457, w36458, w36459, w36460, w36461, w36462, w36463, w36464, w36465, w36466, w36467, w36468, w36469, w36470, w36471, w36472, w36473, w36474, w36475, w36476, w36477, w36478, w36479, w36480, w36481, w36482, w36483, w36484, w36485, w36486, w36487, w36488, w36489, w36490, w36491, w36492, w36493, w36494, w36495, w36496, w36497, w36498, w36499, w36500, w36501, w36502, w36503, w36504, w36505, w36506, w36507, w36508, w36509, w36510, w36511, w36512, w36513, w36514, w36515, w36516, w36517, w36518, w36519, w36520, w36521, w36522, w36523, w36524, w36525, w36526, w36527, w36528, w36529, w36530, w36531, w36532, w36533, w36534, w36535, w36536, w36537, w36538, w36539, w36540, w36541, w36542, w36543, w36544, w36545, w36546, w36547, w36548, w36549, w36550, w36551, w36552, w36553, w36554, w36555, w36556, w36557, w36558, w36559, w36560, w36561, w36562, w36563, w36564, w36565, w36566, w36567, w36568, w36569, w36570, w36571, w36572, w36573, w36574, w36575, w36576, w36577, w36578, w36579, w36580, w36581, w36582, w36583, w36584, w36585, w36586, w36587, w36588, w36589, w36590, w36591, w36592, w36593, w36594, w36595, w36596, w36597, w36598, w36599, w36600, w36601, w36602, w36603, w36604, w36605, w36606, w36607, w36608, w36609, w36610, w36611, w36612, w36613, w36614, w36615, w36616, w36617, w36618, w36619, w36620, w36621, w36622, w36623, w36624, w36625, w36626, w36627, w36628, w36629, w36630, w36631, w36632, w36633, w36634, w36635, w36636, w36637, w36638, w36639, w36640, w36641, w36642, w36643, w36644, w36645, w36646, w36647, w36648, w36649, w36650, w36651, w36652, w36653, w36654, w36655, w36656, w36657, w36658, w36659, w36660, w36661, w36662, w36663, w36664, w36665, w36666, w36667, w36668, w36669, w36670, w36671, w36672, w36673, w36674, w36675, w36676, w36677, w36678, w36679, w36680, w36681, w36682, w36683, w36684, w36685, w36686, w36687, w36688, w36689, w36690, w36691, w36692, w36693, w36694, w36695, w36696, w36697, w36698, w36699, w36700, w36701, w36702, w36703, w36704, w36705, w36706, w36707, w36708, w36709, w36710, w36711, w36712, w36713, w36714, w36715, w36716, w36717, w36718, w36719, w36720, w36721, w36722, w36723, w36724, w36725, w36726, w36727, w36728, w36729, w36730, w36731, w36732, w36733, w36734, w36735, w36736, w36737, w36738, w36739, w36740, w36741, w36742, w36743, w36744, w36745, w36746, w36747, w36748, w36749, w36750, w36751, w36752, w36753, w36754, w36755, w36756, w36757, w36758, w36759, w36760, w36761, w36762, w36763, w36764, w36765, w36766, w36767, w36768, w36769, w36770, w36771, w36772, w36773, w36774, w36775, w36776, w36777, w36778, w36779, w36780, w36781, w36782, w36783, w36784, w36785, w36786, w36787, w36788, w36789, w36790, w36791, w36792, w36793, w36794, w36795, w36796, w36797, w36798, w36799, w36800, w36801, w36802, w36803, w36804, w36805, w36806, w36807, w36808, w36809, w36810, w36811, w36812, w36813, w36814, w36815, w36816, w36817, w36818, w36819, w36820, w36821, w36822, w36823, w36824, w36825, w36826, w36827, w36828, w36829, w36830, w36831, w36832, w36833, w36834, w36835, w36836, w36837, w36838, w36839, w36840, w36841, w36842, w36843, w36844, w36845, w36846, w36847, w36848, w36849, w36850, w36851, w36852, w36853, w36854, w36855, w36856, w36857, w36858, w36859, w36860, w36861, w36862, w36863, w36864, w36865, w36866, w36867, w36868, w36869, w36870, w36871, w36872, w36873, w36874, w36875, w36876, w36877, w36878, w36879, w36880, w36881, w36882, w36883, w36884, w36885, w36886, w36887, w36888, w36889, w36890, w36891, w36892, w36893, w36894, w36895, w36896, w36897, w36898, w36899, w36900, w36901, w36902, w36903, w36904, w36905, w36906, w36907, w36908, w36909, w36910, w36911, w36912, w36913, w36914, w36915, w36916, w36917, w36918, w36919, w36920, w36921, w36922, w36923, w36924, w36925, w36926, w36927, w36928, w36929, w36930, w36931, w36932, w36933, w36934, w36935, w36936, w36937, w36938, w36939, w36940, w36941, w36942, w36943, w36944, w36945, w36946, w36947, w36948, w36949, w36950, w36951, w36952, w36953, w36954, w36955, w36956, w36957, w36958, w36959, w36960, w36961, w36962, w36963, w36964, w36965, w36966, w36967, w36968, w36969, w36970, w36971, w36972, w36973, w36974, w36975, w36976, w36977, w36978, w36979, w36980, w36981, w36982, w36983, w36984, w36985, w36986, w36987, w36988, w36989, w36990, w36991, w36992, w36993, w36994, w36995, w36996, w36997, w36998, w36999, w37000, w37001, w37002, w37003, w37004, w37005, w37006, w37007, w37008, w37009, w37010, w37011, w37012, w37013, w37014, w37015, w37016, w37017, w37018, w37019, w37020, w37021, w37022, w37023, w37024, w37025, w37026, w37027, w37028, w37029, w37030, w37031, w37032, w37033, w37034, w37035, w37036, w37037, w37038, w37039, w37040, w37041, w37042, w37043, w37044, w37045, w37046, w37047, w37048, w37049, w37050, w37051, w37052, w37053, w37054, w37055, w37056, w37057, w37058, w37059, w37060, w37061, w37062, w37063, w37064, w37065, w37066, w37067, w37068, w37069, w37070, w37071, w37072, w37073, w37074, w37075, w37076, w37077, w37078, w37079, w37080, w37081, w37082, w37083, w37084, w37085, w37086, w37087, w37088, w37089, w37090, w37091, w37092, w37093, w37094, w37095, w37096, w37097, w37098, w37099, w37100, w37101, w37102, w37103, w37104, w37105, w37106, w37107, w37108, w37109, w37110, w37111, w37112, w37113, w37114, w37115, w37116, w37117, w37118, w37119, w37120, w37121, w37122, w37123, w37124, w37125, w37126, w37127, w37128, w37129, w37130, w37131, w37132, w37133, w37134, w37135, w37136, w37137, w37138, w37139, w37140, w37141, w37142, w37143, w37144, w37145, w37146, w37147, w37148, w37149, w37150, w37151, w37152, w37153, w37154, w37155, w37156, w37157, w37158, w37159, w37160, w37161, w37162, w37163, w37164, w37165, w37166, w37167, w37168, w37169, w37170, w37171, w37172, w37173, w37174, w37175, w37176, w37177, w37178, w37179, w37180, w37181, w37182, w37183, w37184, w37185, w37186, w37187, w37188, w37189, w37190, w37191, w37192, w37193, w37194, w37195, w37196, w37197, w37198, w37199, w37200, w37201, w37202, w37203, w37204, w37205, w37206, w37207, w37208, w37209, w37210, w37211, w37212, w37213, w37214, w37215, w37216, w37217, w37218, w37219, w37220, w37221, w37222, w37223, w37224, w37225, w37226, w37227, w37228, w37229, w37230, w37231, w37232, w37233, w37234, w37235, w37236, w37237, w37238, w37239, w37240, w37241, w37242, w37243, w37244, w37245, w37246, w37247, w37248, w37249, w37250, w37251, w37252, w37253, w37254, w37255, w37256, w37257, w37258, w37259, w37260, w37261, w37262, w37263, w37264, w37265, w37266, w37267, w37268, w37269, w37270, w37271, w37272, w37273, w37274, w37275, w37276, w37277, w37278, w37279, w37280, w37281, w37282, w37283, w37284, w37285, w37286, w37287, w37288, w37289, w37290, w37291, w37292, w37293, w37294, w37295, w37296, w37297, w37298, w37299, w37300, w37301, w37302, w37303, w37304, w37305, w37306, w37307, w37308, w37309, w37310, w37311, w37312, w37313, w37314, w37315, w37316, w37317, w37318, w37319, w37320, w37321, w37322, w37323, w37324, w37325, w37326, w37327, w37328, w37329, w37330, w37331, w37332, w37333, w37334, w37335, w37336, w37337, w37338, w37339, w37340, w37341, w37342, w37343, w37344, w37345, w37346, w37347, w37348, w37349, w37350, w37351, w37352, w37353, w37354, w37355, w37356, w37357, w37358, w37359, w37360, w37361, w37362, w37363, w37364, w37365, w37366, w37367, w37368, w37369, w37370, w37371, w37372, w37373, w37374, w37375, w37376, w37377, w37378, w37379, w37380, w37381, w37382, w37383, w37384, w37385, w37386, w37387, w37388, w37389, w37390, w37391, w37392, w37393, w37394, w37395, w37396, w37397, w37398, w37399, w37400, w37401, w37402, w37403, w37404, w37405, w37406, w37407, w37408, w37409, w37410, w37411, w37412, w37413, w37414, w37415, w37416, w37417, w37418, w37419, w37420, w37421, w37422, w37423, w37424, w37425, w37426, w37427, w37428, w37429, w37430, w37431, w37432, w37433, w37434, w37435, w37436, w37437, w37438, w37439, w37440, w37441, w37442, w37443, w37444, w37445, w37446, w37447, w37448, w37449, w37450, w37451, w37452, w37453, w37454, w37455, w37456, w37457, w37458, w37459, w37460, w37461, w37462, w37463, w37464, w37465, w37466, w37467, w37468, w37469, w37470, w37471, w37472, w37473, w37474, w37475, w37476, w37477, w37478, w37479, w37480, w37481, w37482, w37483, w37484, w37485, w37486, w37487, w37488, w37489, w37490, w37491, w37492, w37493, w37494, w37495, w37496, w37497, w37498, w37499, w37500, w37501, w37502, w37503, w37504, w37505, w37506, w37507, w37508, w37509, w37510, w37511, w37512, w37513, w37514, w37515, w37516, w37517, w37518, w37519, w37520, w37521, w37522, w37523, w37524, w37525, w37526, w37527, w37528, w37529, w37530, w37531, w37532, w37533, w37534, w37535, w37536, w37537, w37538, w37539, w37540, w37541, w37542, w37543, w37544, w37545, w37546, w37547, w37548, w37549, w37550, w37551, w37552, w37553, w37554, w37555, w37556, w37557, w37558, w37559, w37560, w37561, w37562, w37563, w37564, w37565, w37566, w37567, w37568, w37569, w37570, w37571, w37572, w37573, w37574, w37575, w37576, w37577, w37578, w37579, w37580, w37581, w37582, w37583, w37584, w37585, w37586, w37587, w37588, w37589, w37590, w37591, w37592, w37593, w37594, w37595, w37596, w37597, w37598, w37599, w37600, w37601, w37602, w37603, w37604, w37605, w37606, w37607, w37608, w37609, w37610, w37611, w37612, w37613, w37614, w37615, w37616, w37617, w37618, w37619, w37620, w37621, w37622, w37623, w37624, w37625, w37626, w37627, w37628, w37629, w37630, w37631, w37632, w37633, w37634, w37635, w37636, w37637, w37638, w37639, w37640, w37641, w37642, w37643, w37644, w37645, w37646, w37647, w37648, w37649, w37650, w37651, w37652, w37653, w37654, w37655, w37656, w37657, w37658, w37659, w37660, w37661, w37662, w37663, w37664, w37665, w37666, w37667, w37668, w37669, w37670, w37671, w37672, w37673, w37674, w37675, w37676, w37677, w37678, w37679, w37680, w37681, w37682, w37683, w37684, w37685, w37686, w37687, w37688, w37689, w37690, w37691, w37692, w37693, w37694, w37695, w37696, w37697, w37698, w37699, w37700, w37701, w37702, w37703, w37704, w37705, w37706, w37707, w37708, w37709, w37710, w37711, w37712, w37713, w37714, w37715, w37716, w37717, w37718, w37719, w37720, w37721, w37722, w37723, w37724, w37725, w37726, w37727, w37728, w37729, w37730, w37731, w37732, w37733, w37734, w37735, w37736, w37737, w37738, w37739, w37740, w37741, w37742, w37743, w37744, w37745, w37746, w37747, w37748, w37749, w37750, w37751, w37752, w37753, w37754, w37755, w37756, w37757, w37758, w37759, w37760, w37761, w37762, w37763, w37764, w37765, w37766, w37767, w37768, w37769, w37770, w37771, w37772, w37773, w37774, w37775, w37776, w37777, w37778, w37779, w37780, w37781, w37782, w37783, w37784, w37785, w37786, w37787, w37788, w37789, w37790, w37791, w37792, w37793, w37794, w37795, w37796, w37797, w37798, w37799, w37800, w37801, w37802, w37803, w37804, w37805, w37806, w37807, w37808, w37809, w37810, w37811, w37812, w37813, w37814, w37815, w37816, w37817, w37818, w37819, w37820, w37821, w37822, w37823, w37824, w37825, w37826, w37827, w37828, w37829, w37830, w37831, w37832, w37833, w37834, w37835, w37836, w37837, w37838, w37839, w37840, w37841, w37842, w37843, w37844, w37845, w37846, w37847, w37848, w37849, w37850, w37851, w37852, w37853, w37854, w37855, w37856, w37857, w37858, w37859, w37860, w37861, w37862, w37863, w37864, w37865, w37866, w37867, w37868, w37869, w37870, w37871, w37872, w37873, w37874, w37875, w37876, w37877, w37878, w37879, w37880, w37881, w37882, w37883, w37884, w37885, w37886, w37887, w37888, w37889, w37890, w37891, w37892, w37893, w37894, w37895, w37896, w37897, w37898, w37899, w37900, w37901, w37902, w37903, w37904, w37905, w37906, w37907, w37908, w37909, w37910, w37911, w37912, w37913, w37914, w37915, w37916, w37917, w37918, w37919, w37920, w37921, w37922, w37923, w37924, w37925, w37926, w37927, w37928, w37929, w37930, w37931, w37932, w37933, w37934, w37935, w37936, w37937, w37938, w37939, w37940, w37941, w37942, w37943, w37944, w37945, w37946, w37947, w37948, w37949, w37950, w37951, w37952, w37953, w37954, w37955, w37956, w37957, w37958, w37959, w37960, w37961, w37962, w37963, w37964, w37965, w37966, w37967, w37968, w37969, w37970, w37971, w37972, w37973, w37974, w37975, w37976, w37977, w37978, w37979, w37980, w37981, w37982, w37983, w37984, w37985, w37986, w37987, w37988, w37989, w37990, w37991, w37992, w37993, w37994, w37995, w37996, w37997, w37998, w37999, w38000, w38001, w38002, w38003, w38004, w38005, w38006, w38007, w38008, w38009, w38010, w38011, w38012, w38013, w38014, w38015, w38016, w38017, w38018, w38019, w38020, w38021, w38022, w38023, w38024, w38025, w38026, w38027, w38028, w38029, w38030, w38031, w38032, w38033, w38034, w38035, w38036, w38037, w38038, w38039, w38040, w38041, w38042, w38043, w38044, w38045, w38046, w38047, w38048, w38049, w38050, w38051, w38052, w38053, w38054, w38055, w38056, w38057, w38058, w38059, w38060, w38061, w38062, w38063, w38064, w38065, w38066, w38067, w38068, w38069, w38070, w38071, w38072, w38073, w38074, w38075, w38076, w38077, w38078, w38079, w38080, w38081, w38082, w38083, w38084, w38085, w38086, w38087, w38088, w38089, w38090, w38091, w38092, w38093, w38094, w38095, w38096, w38097, w38098, w38099, w38100, w38101, w38102, w38103, w38104, w38105, w38106, w38107, w38108, w38109, w38110, w38111, w38112, w38113, w38114, w38115, w38116, w38117, w38118, w38119, w38120, w38121, w38122, w38123, w38124, w38125, w38126, w38127, w38128, w38129, w38130, w38131, w38132, w38133, w38134, w38135, w38136, w38137, w38138, w38139, w38140, w38141, w38142, w38143, w38144, w38145, w38146, w38147, w38148, w38149, w38150, w38151, w38152, w38153, w38154, w38155, w38156, w38157, w38158, w38159, w38160, w38161, w38162, w38163, w38164, w38165, w38166, w38167, w38168, w38169, w38170, w38171, w38172, w38173, w38174, w38175, w38176, w38177, w38178, w38179, w38180, w38181, w38182, w38183, w38184, w38185, w38186, w38187, w38188, w38189, w38190, w38191, w38192, w38193, w38194, w38195, w38196, w38197, w38198, w38199, w38200, w38201, w38202, w38203, w38204, w38205, w38206, w38207, w38208, w38209, w38210, w38211, w38212, w38213, w38214, w38215, w38216, w38217, w38218, w38219, w38220, w38221, w38222, w38223, w38224, w38225, w38226, w38227, w38228, w38229, w38230, w38231, w38232, w38233, w38234, w38235, w38236, w38237, w38238, w38239, w38240, w38241, w38242, w38243, w38244, w38245, w38246, w38247, w38248, w38249, w38250, w38251, w38252, w38253, w38254, w38255, w38256, w38257, w38258, w38259, w38260, w38261, w38262, w38263, w38264, w38265, w38266, w38267, w38268, w38269, w38270, w38271, w38272, w38273, w38274, w38275, w38276, w38277, w38278, w38279, w38280, w38281, w38282, w38283, w38284, w38285, w38286, w38287, w38288, w38289, w38290, w38291, w38292, w38293, w38294, w38295, w38296, w38297, w38298, w38299, w38300, w38301, w38302, w38303, w38304, w38305, w38306, w38307, w38308, w38309, w38310, w38311, w38312, w38313, w38314, w38315, w38316, w38317, w38318, w38319, w38320, w38321, w38322, w38323, w38324, w38325, w38326, w38327, w38328, w38329, w38330, w38331, w38332, w38333, w38334, w38335, w38336, w38337, w38338, w38339, w38340, w38341, w38342, w38343, w38344, w38345, w38346, w38347, w38348, w38349, w38350, w38351, w38352, w38353, w38354, w38355, w38356, w38357, w38358, w38359, w38360, w38361, w38362, w38363, w38364, w38365, w38366, w38367, w38368, w38369, w38370, w38371, w38372, w38373, w38374, w38375, w38376, w38377, w38378, w38379, w38380, w38381, w38382, w38383, w38384, w38385, w38386, w38387, w38388, w38389, w38390, w38391, w38392, w38393, w38394, w38395, w38396, w38397, w38398, w38399, w38400, w38401, w38402, w38403, w38404, w38405, w38406, w38407, w38408, w38409, w38410, w38411, w38412, w38413, w38414, w38415, w38416, w38417, w38418, w38419, w38420, w38421, w38422, w38423, w38424, w38425, w38426, w38427, w38428, w38429, w38430, w38431, w38432, w38433, w38434, w38435, w38436, w38437, w38438, w38439, w38440, w38441, w38442, w38443, w38444, w38445, w38446, w38447, w38448, w38449, w38450, w38451, w38452, w38453, w38454, w38455, w38456, w38457, w38458, w38459, w38460, w38461, w38462, w38463, w38464, w38465, w38466, w38467, w38468, w38469, w38470, w38471, w38472, w38473, w38474, w38475, w38476, w38477, w38478, w38479, w38480, w38481, w38482, w38483, w38484, w38485, w38486, w38487, w38488, w38489, w38490, w38491, w38492, w38493, w38494, w38495, w38496, w38497, w38498, w38499, w38500, w38501, w38502, w38503, w38504, w38505, w38506, w38507, w38508, w38509, w38510, w38511, w38512, w38513, w38514, w38515, w38516, w38517, w38518, w38519, w38520, w38521, w38522, w38523, w38524, w38525, w38526, w38527, w38528, w38529, w38530, w38531, w38532, w38533, w38534, w38535, w38536, w38537, w38538, w38539, w38540, w38541, w38542, w38543, w38544, w38545, w38546, w38547, w38548, w38549, w38550, w38551, w38552, w38553, w38554, w38555, w38556, w38557, w38558, w38559, w38560, w38561, w38562, w38563, w38564, w38565, w38566, w38567, w38568, w38569, w38570, w38571, w38572, w38573, w38574, w38575, w38576, w38577, w38578, w38579, w38580, w38581, w38582, w38583, w38584, w38585, w38586, w38587, w38588, w38589, w38590, w38591, w38592, w38593, w38594, w38595, w38596, w38597, w38598, w38599, w38600, w38601, w38602, w38603, w38604, w38605, w38606, w38607, w38608, w38609, w38610, w38611, w38612, w38613, w38614, w38615, w38616, w38617, w38618, w38619, w38620, w38621, w38622, w38623, w38624, w38625, w38626, w38627, w38628, w38629, w38630, w38631, w38632, w38633, w38634, w38635, w38636, w38637, w38638, w38639, w38640, w38641, w38642, w38643, w38644, w38645, w38646, w38647, w38648, w38649, w38650, w38651, w38652, w38653, w38654, w38655, w38656, w38657, w38658, w38659, w38660, w38661, w38662, w38663, w38664, w38665, w38666, w38667, w38668, w38669, w38670, w38671, w38672, w38673, w38674, w38675, w38676, w38677, w38678, w38679, w38680, w38681, w38682, w38683, w38684, w38685, w38686, w38687, w38688, w38689, w38690, w38691, w38692, w38693, w38694, w38695, w38696, w38697, w38698, w38699, w38700, w38701, w38702, w38703, w38704, w38705, w38706, w38707, w38708, w38709, w38710, w38711, w38712, w38713, w38714, w38715, w38716, w38717, w38718, w38719, w38720, w38721, w38722, w38723, w38724, w38725, w38726, w38727, w38728, w38729, w38730, w38731, w38732, w38733, w38734, w38735, w38736, w38737, w38738, w38739, w38740, w38741, w38742, w38743, w38744, w38745, w38746, w38747, w38748, w38749, w38750, w38751, w38752, w38753, w38754, w38755, w38756, w38757, w38758, w38759, w38760, w38761, w38762, w38763, w38764, w38765, w38766, w38767, w38768, w38769, w38770, w38771, w38772, w38773, w38774, w38775, w38776, w38777, w38778, w38779, w38780, w38781, w38782, w38783, w38784, w38785, w38786, w38787, w38788, w38789, w38790, w38791, w38792, w38793, w38794, w38795, w38796, w38797, w38798, w38799, w38800, w38801, w38802, w38803, w38804, w38805, w38806, w38807, w38808, w38809, w38810, w38811, w38812, w38813, w38814, w38815, w38816, w38817, w38818, w38819, w38820, w38821, w38822, w38823, w38824, w38825, w38826, w38827, w38828, w38829, w38830, w38831, w38832, w38833, w38834, w38835, w38836, w38837, w38838, w38839, w38840, w38841, w38842, w38843, w38844, w38845, w38846, w38847, w38848, w38849, w38850, w38851, w38852, w38853, w38854, w38855, w38856, w38857, w38858, w38859, w38860, w38861, w38862, w38863, w38864, w38865, w38866, w38867, w38868, w38869, w38870, w38871, w38872, w38873, w38874, w38875, w38876, w38877, w38878, w38879, w38880, w38881, w38882, w38883, w38884, w38885, w38886, w38887, w38888, w38889, w38890, w38891, w38892, w38893, w38894, w38895, w38896, w38897, w38898, w38899, w38900, w38901, w38902, w38903, w38904, w38905, w38906, w38907, w38908, w38909, w38910, w38911, w38912, w38913, w38914, w38915, w38916, w38917, w38918, w38919, w38920, w38921, w38922, w38923, w38924, w38925, w38926, w38927, w38928, w38929, w38930, w38931, w38932, w38933, w38934, w38935, w38936, w38937, w38938, w38939, w38940, w38941, w38942, w38943, w38944, w38945, w38946, w38947, w38948, w38949, w38950, w38951, w38952, w38953, w38954, w38955, w38956, w38957, w38958, w38959, w38960, w38961, w38962, w38963, w38964, w38965, w38966, w38967, w38968, w38969, w38970, w38971, w38972, w38973, w38974, w38975, w38976, w38977, w38978, w38979, w38980, w38981, w38982, w38983, w38984, w38985, w38986, w38987, w38988, w38989, w38990, w38991, w38992, w38993, w38994, w38995, w38996, w38997, w38998, w38999, w39000, w39001, w39002, w39003, w39004, w39005, w39006, w39007, w39008, w39009, w39010, w39011, w39012, w39013, w39014, w39015, w39016, w39017, w39018, w39019, w39020, w39021, w39022, w39023, w39024, w39025, w39026, w39027, w39028, w39029, w39030, w39031, w39032, w39033, w39034, w39035, w39036, w39037, w39038, w39039, w39040, w39041, w39042, w39043, w39044, w39045, w39046, w39047, w39048, w39049, w39050, w39051, w39052, w39053, w39054, w39055, w39056, w39057, w39058, w39059, w39060, w39061, w39062, w39063, w39064, w39065, w39066, w39067, w39068, w39069, w39070, w39071, w39072, w39073, w39074, w39075, w39076, w39077, w39078, w39079, w39080, w39081, w39082, w39083, w39084, w39085, w39086, w39087, w39088, w39089, w39090, w39091, w39092, w39093, w39094, w39095, w39096, w39097, w39098, w39099, w39100, w39101, w39102, w39103, w39104, w39105, w39106, w39107, w39108, w39109, w39110, w39111, w39112, w39113, w39114, w39115, w39116, w39117, w39118, w39119, w39120, w39121, w39122, w39123, w39124, w39125, w39126, w39127, w39128, w39129, w39130, w39131, w39132, w39133, w39134, w39135, w39136, w39137, w39138, w39139, w39140, w39141, w39142, w39143, w39144, w39145, w39146, w39147, w39148, w39149, w39150, w39151, w39152, w39153, w39154, w39155, w39156, w39157, w39158, w39159, w39160, w39161, w39162, w39163, w39164, w39165, w39166, w39167, w39168, w39169, w39170, w39171, w39172, w39173, w39174, w39175, w39176, w39177, w39178, w39179, w39180, w39181, w39182, w39183, w39184, w39185, w39186, w39187, w39188, w39189, w39190, w39191, w39192, w39193, w39194, w39195, w39196, w39197, w39198, w39199, w39200, w39201, w39202, w39203, w39204, w39205, w39206, w39207, w39208, w39209, w39210, w39211, w39212, w39213, w39214, w39215, w39216, w39217, w39218, w39219, w39220, w39221, w39222, w39223, w39224, w39225, w39226, w39227, w39228, w39229, w39230, w39231, w39232, w39233, w39234, w39235, w39236, w39237, w39238, w39239, w39240, w39241, w39242, w39243, w39244, w39245, w39246, w39247, w39248, w39249, w39250, w39251, w39252, w39253, w39254, w39255, w39256, w39257, w39258, w39259, w39260, w39261, w39262, w39263, w39264, w39265, w39266, w39267, w39268, w39269, w39270, w39271, w39272, w39273, w39274, w39275, w39276, w39277, w39278, w39279, w39280, w39281, w39282, w39283, w39284, w39285, w39286, w39287, w39288, w39289, w39290, w39291, w39292, w39293, w39294, w39295, w39296, w39297, w39298, w39299, w39300, w39301, w39302, w39303, w39304, w39305, w39306, w39307, w39308, w39309, w39310, w39311, w39312, w39313, w39314, w39315, w39316, w39317, w39318, w39319, w39320, w39321, w39322, w39323, w39324, w39325, w39326, w39327, w39328, w39329, w39330, w39331, w39332, w39333, w39334, w39335, w39336, w39337, w39338, w39339, w39340, w39341, w39342, w39343, w39344, w39345, w39346, w39347, w39348, w39349, w39350, w39351, w39352, w39353, w39354, w39355, w39356, w39357, w39358, w39359, w39360, w39361, w39362, w39363, w39364, w39365, w39366, w39367, w39368, w39369, w39370, w39371, w39372, w39373, w39374, w39375, w39376, w39377, w39378, w39379, w39380, w39381, w39382, w39383, w39384, w39385, w39386, w39387, w39388, w39389, w39390, w39391, w39392, w39393, w39394, w39395, w39396, w39397, w39398, w39399, w39400, w39401, w39402, w39403, w39404, w39405, w39406, w39407, w39408, w39409, w39410, w39411, w39412, w39413, w39414, w39415, w39416, w39417, w39418, w39419, w39420, w39421, w39422, w39423, w39424, w39425, w39426, w39427, w39428, w39429, w39430, w39431, w39432, w39433, w39434, w39435, w39436, w39437, w39438, w39439, w39440, w39441, w39442, w39443, w39444, w39445, w39446, w39447, w39448, w39449, w39450, w39451, w39452, w39453, w39454, w39455, w39456, w39457, w39458, w39459, w39460, w39461, w39462, w39463, w39464, w39465, w39466, w39467, w39468, w39469, w39470, w39471, w39472, w39473, w39474, w39475, w39476, w39477, w39478, w39479, w39480, w39481, w39482, w39483, w39484, w39485, w39486, w39487, w39488, w39489, w39490, w39491, w39492, w39493, w39494, w39495, w39496, w39497, w39498, w39499, w39500, w39501, w39502, w39503, w39504, w39505, w39506, w39507, w39508, w39509, w39510, w39511, w39512, w39513, w39514, w39515, w39516, w39517, w39518, w39519, w39520, w39521, w39522, w39523, w39524, w39525, w39526, w39527, w39528, w39529, w39530, w39531, w39532, w39533, w39534, w39535, w39536, w39537, w39538, w39539, w39540, w39541, w39542, w39543, w39544, w39545, w39546, w39547, w39548, w39549, w39550, w39551, w39552, w39553, w39554, w39555, w39556, w39557, w39558, w39559, w39560, w39561, w39562, w39563, w39564, w39565, w39566, w39567, w39568, w39569, w39570, w39571, w39572, w39573, w39574, w39575, w39576, w39577, w39578, w39579, w39580, w39581, w39582, w39583, w39584, w39585, w39586, w39587, w39588, w39589, w39590, w39591, w39592, w39593, w39594, w39595, w39596, w39597, w39598, w39599, w39600, w39601, w39602, w39603, w39604, w39605, w39606, w39607, w39608, w39609, w39610, w39611, w39612, w39613, w39614, w39615, w39616, w39617, w39618, w39619, w39620, w39621, w39622, w39623, w39624, w39625, w39626, w39627, w39628, w39629, w39630, w39631, w39632, w39633, w39634, w39635, w39636, w39637, w39638, w39639, w39640, w39641, w39642, w39643, w39644, w39645, w39646, w39647, w39648, w39649, w39650, w39651, w39652, w39653, w39654, w39655, w39656, w39657, w39658, w39659, w39660, w39661, w39662, w39663, w39664, w39665, w39666, w39667, w39668, w39669, w39670, w39671, w39672, w39673, w39674, w39675, w39676, w39677, w39678, w39679, w39680, w39681, w39682, w39683, w39684, w39685, w39686, w39687, w39688, w39689, w39690, w39691, w39692, w39693, w39694, w39695, w39696, w39697, w39698, w39699, w39700, w39701, w39702, w39703, w39704, w39705, w39706, w39707, w39708, w39709, w39710, w39711, w39712, w39713, w39714, w39715, w39716, w39717, w39718, w39719, w39720, w39721, w39722, w39723, w39724, w39725, w39726, w39727, w39728, w39729, w39730, w39731, w39732, w39733, w39734, w39735, w39736, w39737, w39738, w39739, w39740, w39741, w39742, w39743, w39744, w39745, w39746, w39747, w39748, w39749, w39750, w39751, w39752, w39753, w39754, w39755, w39756, w39757, w39758, w39759, w39760, w39761, w39762, w39763, w39764, w39765, w39766, w39767, w39768, w39769, w39770, w39771, w39772, w39773, w39774, w39775, w39776, w39777, w39778, w39779, w39780, w39781, w39782, w39783, w39784, w39785, w39786, w39787, w39788, w39789, w39790, w39791, w39792, w39793, w39794, w39795, w39796, w39797, w39798, w39799, w39800, w39801, w39802, w39803, w39804, w39805, w39806, w39807, w39808, w39809, w39810, w39811, w39812, w39813, w39814, w39815, w39816, w39817, w39818, w39819, w39820, w39821, w39822, w39823, w39824, w39825, w39826, w39827, w39828, w39829, w39830, w39831, w39832, w39833, w39834, w39835, w39836, w39837, w39838, w39839, w39840, w39841, w39842, w39843, w39844, w39845, w39846, w39847, w39848, w39849, w39850, w39851, w39852, w39853, w39854, w39855, w39856, w39857, w39858, w39859, w39860, w39861, w39862, w39863, w39864, w39865, w39866, w39867, w39868, w39869, w39870, w39871, w39872, w39873, w39874, w39875, w39876, w39877, w39878, w39879, w39880, w39881, w39882, w39883, w39884, w39885, w39886, w39887, w39888, w39889, w39890, w39891, w39892, w39893, w39894, w39895, w39896, w39897, w39898, w39899, w39900, w39901, w39902, w39903, w39904, w39905, w39906, w39907, w39908, w39909, w39910, w39911, w39912, w39913, w39914, w39915, w39916, w39917, w39918, w39919, w39920, w39921, w39922, w39923, w39924, w39925, w39926, w39927, w39928, w39929, w39930, w39931, w39932, w39933, w39934, w39935, w39936, w39937, w39938, w39939, w39940, w39941, w39942, w39943, w39944, w39945, w39946, w39947, w39948, w39949, w39950, w39951, w39952, w39953, w39954, w39955, w39956, w39957, w39958, w39959, w39960, w39961, w39962, w39963, w39964, w39965, w39966, w39967, w39968, w39969, w39970, w39971, w39972, w39973, w39974, w39975, w39976, w39977, w39978, w39979, w39980, w39981, w39982, w39983, w39984, w39985, w39986, w39987, w39988, w39989, w39990, w39991, w39992, w39993, w39994, w39995, w39996, w39997, w39998, w39999, w40000, w40001, w40002, w40003, w40004, w40005, w40006, w40007, w40008, w40009, w40010, w40011, w40012, w40013, w40014, w40015, w40016, w40017, w40018, w40019, w40020, w40021, w40022, w40023, w40024, w40025, w40026, w40027, w40028, w40029, w40030, w40031, w40032, w40033, w40034, w40035, w40036, w40037, w40038, w40039, w40040, w40041, w40042, w40043, w40044, w40045, w40046, w40047, w40048, w40049, w40050, w40051, w40052, w40053, w40054, w40055, w40056, w40057, w40058, w40059, w40060, w40061, w40062, w40063, w40064, w40065, w40066, w40067, w40068, w40069, w40070, w40071, w40072, w40073, w40074, w40075, w40076, w40077, w40078, w40079, w40080, w40081, w40082, w40083, w40084, w40085, w40086, w40087, w40088, w40089, w40090, w40091, w40092, w40093, w40094, w40095, w40096, w40097, w40098, w40099, w40100, w40101, w40102, w40103, w40104, w40105, w40106, w40107, w40108, w40109, w40110, w40111, w40112, w40113, w40114, w40115, w40116, w40117, w40118, w40119, w40120, w40121, w40122, w40123, w40124, w40125, w40126, w40127, w40128, w40129, w40130, w40131, w40132, w40133, w40134, w40135, w40136, w40137, w40138, w40139, w40140, w40141, w40142, w40143, w40144, w40145, w40146, w40147, w40148, w40149, w40150, w40151, w40152, w40153, w40154, w40155, w40156, w40157, w40158, w40159, w40160, w40161, w40162, w40163, w40164, w40165, w40166, w40167, w40168, w40169, w40170, w40171, w40172, w40173, w40174, w40175, w40176, w40177, w40178, w40179, w40180, w40181, w40182, w40183, w40184, w40185, w40186, w40187, w40188, w40189, w40190, w40191, w40192, w40193, w40194, w40195, w40196, w40197, w40198, w40199, w40200, w40201, w40202, w40203, w40204, w40205, w40206, w40207, w40208, w40209, w40210, w40211, w40212, w40213, w40214, w40215, w40216, w40217, w40218, w40219, w40220, w40221, w40222, w40223, w40224, w40225, w40226, w40227, w40228, w40229, w40230, w40231, w40232, w40233, w40234, w40235, w40236, w40237, w40238, w40239, w40240, w40241, w40242, w40243, w40244, w40245, w40246, w40247, w40248, w40249, w40250, w40251, w40252, w40253, w40254, w40255, w40256, w40257, w40258, w40259, w40260, w40261, w40262, w40263, w40264, w40265, w40266, w40267, w40268, w40269, w40270, w40271, w40272, w40273, w40274, w40275, w40276, w40277, w40278, w40279, w40280, w40281, w40282, w40283, w40284, w40285, w40286, w40287, w40288, w40289, w40290, w40291, w40292, w40293, w40294, w40295, w40296, w40297, w40298, w40299, w40300, w40301, w40302, w40303, w40304, w40305, w40306, w40307, w40308, w40309, w40310, w40311, w40312, w40313, w40314, w40315, w40316, w40317, w40318, w40319, w40320, w40321, w40322, w40323, w40324, w40325, w40326, w40327, w40328, w40329, w40330, w40331, w40332, w40333, w40334, w40335, w40336, w40337, w40338, w40339, w40340, w40341, w40342, w40343, w40344, w40345, w40346, w40347, w40348, w40349, w40350, w40351, w40352, w40353, w40354, w40355, w40356, w40357, w40358, w40359, w40360, w40361, w40362, w40363, w40364, w40365, w40366, w40367, w40368, w40369, w40370, w40371, w40372, w40373, w40374, w40375, w40376, w40377, w40378, w40379, w40380, w40381, w40382, w40383, w40384, w40385, w40386, w40387, w40388, w40389, w40390, w40391, w40392, w40393, w40394, w40395, w40396, w40397, w40398, w40399, w40400, w40401, w40402, w40403, w40404, w40405, w40406, w40407, w40408, w40409, w40410, w40411, w40412, w40413, w40414, w40415, w40416, w40417, w40418, w40419, w40420, w40421, w40422, w40423, w40424, w40425, w40426, w40427, w40428, w40429, w40430, w40431, w40432, w40433, w40434, w40435, w40436, w40437, w40438, w40439, w40440, w40441, w40442, w40443, w40444, w40445, w40446, w40447, w40448, w40449, w40450, w40451, w40452, w40453, w40454, w40455, w40456, w40457, w40458, w40459, w40460, w40461, w40462, w40463, w40464, w40465, w40466, w40467, w40468, w40469, w40470, w40471, w40472, w40473, w40474, w40475, w40476, w40477, w40478, w40479, w40480, w40481, w40482, w40483, w40484, w40485, w40486, w40487, w40488, w40489, w40490, w40491, w40492, w40493, w40494, w40495, w40496, w40497, w40498, w40499, w40500, w40501, w40502, w40503, w40504, w40505, w40506, w40507, w40508, w40509, w40510, w40511, w40512, w40513, w40514, w40515, w40516, w40517, w40518, w40519, w40520, w40521, w40522, w40523, w40524, w40525, w40526, w40527, w40528, w40529, w40530, w40531, w40532, w40533, w40534, w40535, w40536, w40537, w40538, w40539, w40540, w40541, w40542, w40543, w40544, w40545, w40546, w40547, w40548, w40549, w40550, w40551, w40552, w40553, w40554, w40555, w40556, w40557, w40558, w40559, w40560, w40561, w40562, w40563, w40564, w40565, w40566, w40567, w40568, w40569, w40570, w40571, w40572, w40573, w40574, w40575, w40576, w40577, w40578, w40579, w40580, w40581, w40582, w40583, w40584, w40585, w40586, w40587, w40588, w40589, w40590, w40591, w40592, w40593, w40594, w40595, w40596, w40597, w40598, w40599, w40600, w40601, w40602, w40603, w40604, w40605, w40606, w40607, w40608, w40609, w40610, w40611, w40612, w40613, w40614, w40615, w40616, w40617, w40618, w40619, w40620, w40621, w40622, w40623, w40624, w40625, w40626, w40627, w40628, w40629, w40630, w40631, w40632, w40633, w40634, w40635, w40636, w40637, w40638, w40639, w40640, w40641, w40642, w40643, w40644, w40645, w40646, w40647, w40648, w40649, w40650, w40651, w40652, w40653, w40654, w40655, w40656, w40657, w40658, w40659, w40660, w40661, w40662, w40663, w40664, w40665, w40666, w40667, w40668, w40669, w40670, w40671, w40672, w40673, w40674, w40675, w40676, w40677, w40678, w40679, w40680, w40681, w40682, w40683, w40684, w40685, w40686, w40687, w40688, w40689, w40690, w40691, w40692, w40693, w40694, w40695, w40696, w40697, w40698, w40699, w40700, w40701, w40702, w40703, w40704, w40705, w40706, w40707, w40708, w40709, w40710, w40711, w40712, w40713, w40714, w40715, w40716, w40717, w40718, w40719, w40720, w40721, w40722, w40723, w40724, w40725, w40726, w40727, w40728, w40729, w40730, w40731, w40732, w40733, w40734, w40735, w40736, w40737, w40738, w40739, w40740, w40741, w40742, w40743, w40744, w40745, w40746, w40747, w40748, w40749, w40750, w40751, w40752, w40753, w40754, w40755, w40756, w40757, w40758, w40759, w40760, w40761, w40762, w40763, w40764, w40765, w40766, w40767, w40768, w40769, w40770, w40771, w40772, w40773, w40774, w40775, w40776, w40777, w40778, w40779, w40780, w40781, w40782, w40783, w40784, w40785, w40786, w40787, w40788, w40789, w40790, w40791, w40792, w40793, w40794, w40795, w40796, w40797, w40798, w40799, w40800, w40801, w40802, w40803, w40804, w40805, w40806, w40807, w40808, w40809, w40810, w40811, w40812, w40813, w40814, w40815, w40816, w40817, w40818, w40819, w40820, w40821, w40822, w40823, w40824, w40825, w40826, w40827, w40828, w40829, w40830, w40831, w40832, w40833, w40834, w40835, w40836, w40837, w40838, w40839, w40840, w40841, w40842, w40843, w40844, w40845, w40846, w40847, w40848, w40849, w40850, w40851, w40852, w40853, w40854, w40855, w40856, w40857, w40858, w40859, w40860, w40861, w40862, w40863, w40864, w40865, w40866, w40867, w40868, w40869, w40870, w40871, w40872, w40873, w40874, w40875, w40876, w40877, w40878, w40879, w40880, w40881, w40882, w40883, w40884, w40885, w40886, w40887, w40888, w40889, w40890, w40891, w40892, w40893, w40894, w40895, w40896, w40897, w40898, w40899, w40900, w40901, w40902, w40903, w40904, w40905, w40906, w40907, w40908, w40909, w40910, w40911, w40912, w40913, w40914, w40915, w40916, w40917, w40918, w40919, w40920, w40921, w40922, w40923, w40924, w40925, w40926, w40927, w40928, w40929, w40930, w40931, w40932, w40933, w40934, w40935, w40936, w40937, w40938, w40939, w40940, w40941, w40942, w40943, w40944, w40945, w40946, w40947, w40948, w40949, w40950, w40951, w40952, w40953, w40954, w40955, w40956, w40957, w40958, w40959, w40960, w40961, w40962, w40963, w40964, w40965, w40966, w40967, w40968, w40969, w40970, w40971, w40972, w40973, w40974, w40975, w40976, w40977, w40978, w40979, w40980, w40981, w40982, w40983, w40984, w40985, w40986, w40987, w40988, w40989, w40990, w40991, w40992, w40993, w40994, w40995, w40996, w40997, w40998, w40999, w41000, w41001, w41002, w41003, w41004, w41005, w41006, w41007, w41008, w41009, w41010, w41011, w41012, w41013, w41014, w41015, w41016, w41017, w41018, w41019, w41020, w41021, w41022, w41023, w41024, w41025, w41026, w41027, w41028, w41029, w41030, w41031, w41032, w41033, w41034, w41035, w41036, w41037, w41038, w41039, w41040, w41041, w41042, w41043, w41044, w41045, w41046, w41047, w41048, w41049, w41050, w41051, w41052, w41053, w41054, w41055, w41056, w41057, w41058, w41059, w41060, w41061, w41062, w41063, w41064, w41065, w41066, w41067, w41068, w41069, w41070, w41071, w41072, w41073, w41074, w41075, w41076, w41077, w41078, w41079, w41080, w41081, w41082, w41083, w41084, w41085, w41086, w41087, w41088, w41089, w41090, w41091, w41092, w41093, w41094, w41095, w41096, w41097, w41098, w41099, w41100, w41101, w41102, w41103, w41104, w41105, w41106, w41107, w41108, w41109, w41110, w41111, w41112, w41113, w41114, w41115, w41116, w41117, w41118, w41119, w41120, w41121, w41122, w41123, w41124, w41125, w41126, w41127, w41128, w41129, w41130, w41131, w41132, w41133, w41134, w41135, w41136, w41137, w41138, w41139, w41140, w41141, w41142, w41143, w41144, w41145, w41146, w41147, w41148, w41149, w41150, w41151, w41152, w41153, w41154, w41155, w41156, w41157, w41158, w41159, w41160, w41161, w41162, w41163, w41164, w41165, w41166, w41167, w41168, w41169, w41170, w41171, w41172, w41173, w41174, w41175, w41176, w41177, w41178, w41179, w41180, w41181, w41182, w41183, w41184, w41185, w41186, w41187, w41188, w41189, w41190, w41191, w41192, w41193, w41194, w41195, w41196, w41197, w41198, w41199, w41200, w41201, w41202, w41203, w41204, w41205, w41206, w41207, w41208, w41209, w41210, w41211, w41212, w41213, w41214, w41215, w41216, w41217, w41218, w41219, w41220, w41221, w41222, w41223, w41224, w41225, w41226, w41227, w41228, w41229, w41230, w41231, w41232, w41233, w41234, w41235, w41236, w41237, w41238, w41239, w41240, w41241, w41242, w41243, w41244, w41245, w41246, w41247, w41248, w41249, w41250, w41251, w41252, w41253, w41254, w41255, w41256, w41257, w41258, w41259, w41260, w41261, w41262, w41263, w41264, w41265, w41266, w41267, w41268, w41269, w41270, w41271, w41272, w41273, w41274, w41275, w41276, w41277, w41278, w41279, w41280, w41281, w41282, w41283, w41284, w41285, w41286, w41287, w41288, w41289, w41290, w41291, w41292, w41293, w41294, w41295, w41296, w41297, w41298, w41299, w41300, w41301, w41302, w41303, w41304, w41305, w41306, w41307, w41308, w41309, w41310, w41311, w41312, w41313, w41314, w41315, w41316, w41317, w41318, w41319, w41320, w41321, w41322, w41323, w41324, w41325, w41326, w41327, w41328, w41329, w41330, w41331, w41332, w41333, w41334, w41335, w41336, w41337, w41338, w41339, w41340, w41341, w41342, w41343, w41344, w41345, w41346, w41347, w41348, w41349, w41350, w41351, w41352, w41353, w41354, w41355, w41356, w41357, w41358, w41359, w41360, w41361, w41362, w41363, w41364, w41365, w41366, w41367, w41368, w41369, w41370, w41371, w41372, w41373, w41374, w41375, w41376, w41377, w41378, w41379, w41380, w41381, w41382, w41383, w41384, w41385, w41386, w41387, w41388, w41389, w41390, w41391, w41392, w41393, w41394, w41395, w41396, w41397, w41398, w41399, w41400, w41401, w41402, w41403, w41404, w41405, w41406, w41407, w41408, w41409, w41410, w41411, w41412, w41413, w41414, w41415, w41416, w41417, w41418, w41419, w41420, w41421, w41422, w41423, w41424, w41425, w41426, w41427, w41428, w41429, w41430, w41431, w41432, w41433, w41434, w41435, w41436, w41437, w41438, w41439, w41440, w41441, w41442, w41443, w41444, w41445, w41446, w41447, w41448, w41449, w41450, w41451, w41452, w41453, w41454, w41455, w41456, w41457, w41458, w41459, w41460, w41461, w41462, w41463, w41464, w41465, w41466, w41467, w41468, w41469, w41470, w41471, w41472, w41473, w41474, w41475, w41476, w41477, w41478, w41479, w41480, w41481, w41482, w41483, w41484, w41485, w41486, w41487, w41488, w41489, w41490, w41491, w41492, w41493, w41494, w41495, w41496, w41497, w41498, w41499, w41500, w41501, w41502, w41503, w41504, w41505, w41506, w41507, w41508, w41509, w41510, w41511, w41512, w41513, w41514, w41515, w41516, w41517, w41518, w41519, w41520, w41521, w41522, w41523, w41524, w41525, w41526, w41527, w41528, w41529, w41530, w41531, w41532, w41533, w41534, w41535, w41536, w41537, w41538, w41539, w41540, w41541, w41542, w41543, w41544, w41545, w41546, w41547, w41548, w41549, w41550, w41551, w41552, w41553, w41554, w41555, w41556, w41557, w41558, w41559, w41560, w41561, w41562, w41563, w41564, w41565, w41566, w41567, w41568, w41569, w41570, w41571, w41572, w41573, w41574, w41575, w41576, w41577, w41578, w41579, w41580, w41581, w41582, w41583, w41584, w41585, w41586, w41587, w41588, w41589, w41590, w41591, w41592, w41593, w41594, w41595, w41596, w41597, w41598, w41599, w41600, w41601, w41602, w41603, w41604, w41605, w41606, w41607, w41608, w41609, w41610, w41611, w41612, w41613, w41614, w41615, w41616, w41617, w41618, w41619, w41620, w41621, w41622, w41623, w41624, w41625, w41626, w41627, w41628, w41629, w41630, w41631, w41632, w41633, w41634, w41635, w41636, w41637, w41638, w41639, w41640, w41641, w41642, w41643, w41644, w41645, w41646, w41647, w41648, w41649, w41650, w41651, w41652, w41653, w41654, w41655, w41656, w41657, w41658, w41659, w41660, w41661, w41662, w41663, w41664, w41665, w41666, w41667, w41668, w41669, w41670, w41671, w41672, w41673, w41674, w41675, w41676, w41677, w41678, w41679, w41680, w41681, w41682, w41683, w41684, w41685, w41686, w41687, w41688, w41689, w41690, w41691, w41692, w41693, w41694, w41695, w41696, w41697, w41698, w41699, w41700, w41701, w41702, w41703, w41704, w41705, w41706, w41707, w41708, w41709, w41710, w41711, w41712, w41713, w41714, w41715, w41716, w41717, w41718, w41719, w41720, w41721, w41722, w41723, w41724, w41725, w41726, w41727, w41728, w41729, w41730, w41731, w41732, w41733, w41734, w41735, w41736, w41737, w41738, w41739, w41740, w41741, w41742, w41743, w41744, w41745, w41746, w41747, w41748, w41749, w41750, w41751, w41752, w41753, w41754, w41755, w41756, w41757, w41758, w41759, w41760, w41761, w41762, w41763, w41764, w41765, w41766, w41767, w41768, w41769, w41770, w41771, w41772, w41773, w41774, w41775, w41776, w41777, w41778, w41779, w41780, w41781, w41782, w41783, w41784, w41785, w41786, w41787, w41788, w41789, w41790, w41791, w41792, w41793, w41794, w41795, w41796, w41797, w41798, w41799, w41800, w41801, w41802, w41803, w41804, w41805, w41806, w41807, w41808, w41809, w41810, w41811, w41812, w41813, w41814, w41815, w41816, w41817, w41818, w41819, w41820, w41821, w41822, w41823, w41824, w41825, w41826, w41827, w41828, w41829, w41830, w41831, w41832, w41833, w41834, w41835, w41836, w41837, w41838, w41839, w41840, w41841, w41842, w41843, w41844, w41845, w41846, w41847, w41848, w41849, w41850, w41851, w41852, w41853, w41854, w41855, w41856, w41857, w41858, w41859, w41860, w41861, w41862, w41863, w41864, w41865, w41866, w41867, w41868, w41869, w41870, w41871, w41872, w41873, w41874, w41875, w41876, w41877, w41878, w41879, w41880, w41881, w41882, w41883, w41884, w41885, w41886, w41887, w41888, w41889, w41890, w41891, w41892, w41893, w41894, w41895, w41896, w41897, w41898, w41899, w41900, w41901, w41902, w41903, w41904, w41905, w41906, w41907, w41908, w41909, w41910, w41911, w41912, w41913, w41914, w41915, w41916, w41917, w41918, w41919, w41920, w41921, w41922, w41923, w41924, w41925, w41926, w41927, w41928, w41929, w41930, w41931, w41932, w41933, w41934, w41935, w41936, w41937, w41938, w41939, w41940, w41941, w41942, w41943, w41944, w41945, w41946, w41947, w41948, w41949, w41950, w41951, w41952, w41953, w41954, w41955, w41956, w41957, w41958, w41959, w41960, w41961, w41962, w41963, w41964, w41965, w41966, w41967, w41968, w41969, w41970, w41971, w41972, w41973, w41974, w41975, w41976, w41977, w41978, w41979, w41980, w41981, w41982, w41983, w41984, w41985, w41986, w41987, w41988, w41989, w41990, w41991, w41992, w41993, w41994, w41995, w41996, w41997, w41998, w41999, w42000, w42001, w42002, w42003, w42004, w42005, w42006, w42007, w42008, w42009, w42010, w42011, w42012, w42013, w42014, w42015, w42016, w42017, w42018, w42019, w42020, w42021, w42022, w42023, w42024, w42025, w42026, w42027, w42028, w42029, w42030, w42031, w42032, w42033, w42034, w42035, w42036, w42037, w42038, w42039, w42040, w42041, w42042, w42043, w42044, w42045, w42046, w42047, w42048, w42049, w42050, w42051, w42052, w42053, w42054, w42055, w42056, w42057, w42058, w42059, w42060, w42061, w42062, w42063, w42064, w42065, w42066, w42067, w42068, w42069, w42070, w42071, w42072, w42073, w42074, w42075, w42076, w42077, w42078, w42079, w42080, w42081, w42082, w42083, w42084, w42085, w42086, w42087, w42088, w42089, w42090, w42091, w42092, w42093, w42094, w42095, w42096, w42097, w42098, w42099, w42100, w42101, w42102, w42103, w42104, w42105, w42106, w42107, w42108, w42109, w42110, w42111, w42112, w42113, w42114, w42115, w42116, w42117, w42118, w42119, w42120, w42121, w42122, w42123, w42124, w42125, w42126, w42127, w42128, w42129, w42130, w42131, w42132, w42133, w42134, w42135, w42136, w42137, w42138, w42139, w42140, w42141, w42142, w42143, w42144, w42145, w42146, w42147, w42148, w42149, w42150, w42151, w42152, w42153, w42154, w42155, w42156, w42157, w42158, w42159, w42160, w42161, w42162, w42163, w42164, w42165, w42166, w42167, w42168, w42169, w42170, w42171, w42172, w42173, w42174, w42175, w42176, w42177, w42178, w42179, w42180, w42181, w42182, w42183, w42184, w42185, w42186, w42187, w42188, w42189, w42190, w42191, w42192, w42193, w42194, w42195, w42196, w42197, w42198, w42199, w42200, w42201, w42202, w42203, w42204, w42205, w42206, w42207, w42208, w42209, w42210, w42211, w42212, w42213, w42214, w42215, w42216, w42217, w42218, w42219, w42220, w42221, w42222, w42223, w42224, w42225, w42226, w42227, w42228, w42229, w42230, w42231, w42232, w42233, w42234, w42235, w42236, w42237, w42238, w42239, w42240, w42241, w42242, w42243, w42244, w42245, w42246, w42247, w42248, w42249, w42250, w42251, w42252, w42253, w42254, w42255, w42256, w42257, w42258, w42259, w42260, w42261, w42262, w42263, w42264, w42265, w42266, w42267, w42268, w42269, w42270, w42271, w42272, w42273, w42274, w42275, w42276, w42277, w42278, w42279, w42280, w42281, w42282, w42283, w42284, w42285, w42286, w42287, w42288, w42289, w42290, w42291, w42292, w42293, w42294, w42295, w42296, w42297, w42298, w42299, w42300, w42301, w42302, w42303, w42304, w42305, w42306, w42307, w42308, w42309, w42310, w42311, w42312, w42313, w42314, w42315, w42316, w42317, w42318, w42319, w42320, w42321, w42322, w42323, w42324, w42325, w42326, w42327, w42328, w42329, w42330, w42331, w42332, w42333, w42334, w42335, w42336, w42337, w42338, w42339, w42340, w42341, w42342, w42343, w42344, w42345, w42346, w42347, w42348, w42349, w42350, w42351, w42352, w42353, w42354, w42355, w42356, w42357, w42358, w42359, w42360, w42361, w42362, w42363, w42364, w42365, w42366, w42367, w42368, w42369, w42370, w42371, w42372, w42373, w42374, w42375, w42376, w42377, w42378, w42379, w42380, w42381, w42382, w42383, w42384, w42385, w42386, w42387, w42388, w42389, w42390, w42391, w42392, w42393, w42394, w42395, w42396, w42397, w42398, w42399, w42400, w42401, w42402, w42403, w42404, w42405, w42406, w42407, w42408, w42409, w42410, w42411, w42412, w42413, w42414, w42415, w42416, w42417, w42418, w42419, w42420, w42421, w42422, w42423, w42424, w42425, w42426, w42427, w42428, w42429, w42430, w42431, w42432, w42433, w42434, w42435, w42436, w42437, w42438, w42439, w42440, w42441, w42442, w42443, w42444, w42445, w42446, w42447, w42448, w42449, w42450, w42451, w42452, w42453, w42454, w42455, w42456, w42457, w42458, w42459, w42460, w42461, w42462, w42463, w42464, w42465, w42466, w42467, w42468, w42469, w42470, w42471, w42472, w42473, w42474, w42475, w42476, w42477, w42478, w42479, w42480, w42481, w42482, w42483, w42484, w42485, w42486, w42487, w42488, w42489, w42490, w42491, w42492, w42493, w42494, w42495, w42496, w42497, w42498, w42499, w42500, w42501, w42502, w42503, w42504, w42505, w42506, w42507, w42508, w42509, w42510, w42511, w42512, w42513, w42514, w42515, w42516, w42517, w42518, w42519, w42520, w42521, w42522, w42523, w42524, w42525, w42526, w42527, w42528, w42529, w42530, w42531, w42532, w42533, w42534, w42535, w42536, w42537, w42538, w42539, w42540, w42541, w42542, w42543, w42544, w42545, w42546, w42547, w42548, w42549, w42550, w42551, w42552, w42553, w42554, w42555, w42556, w42557, w42558, w42559, w42560, w42561, w42562, w42563, w42564, w42565, w42566, w42567, w42568, w42569, w42570, w42571, w42572, w42573, w42574, w42575, w42576, w42577, w42578, w42579, w42580, w42581, w42582, w42583, w42584, w42585, w42586, w42587, w42588, w42589, w42590, w42591, w42592, w42593, w42594, w42595, w42596, w42597, w42598, w42599, w42600, w42601, w42602, w42603, w42604, w42605, w42606, w42607, w42608, w42609, w42610, w42611, w42612, w42613, w42614, w42615, w42616, w42617, w42618, w42619, w42620, w42621, w42622, w42623, w42624, w42625, w42626, w42627, w42628, w42629, w42630, w42631, w42632, w42633, w42634, w42635, w42636, w42637, w42638, w42639, w42640, w42641, w42642, w42643, w42644, w42645, w42646, w42647, w42648, w42649, w42650, w42651, w42652, w42653, w42654, w42655, w42656, w42657, w42658, w42659, w42660, w42661, w42662, w42663, w42664, w42665, w42666, w42667, w42668, w42669, w42670, w42671, w42672, w42673, w42674, w42675, w42676, w42677, w42678, w42679, w42680, w42681, w42682, w42683, w42684, w42685, w42686, w42687, w42688, w42689, w42690, w42691, w42692, w42693, w42694, w42695, w42696, w42697, w42698, w42699, w42700, w42701, w42702, w42703, w42704, w42705, w42706, w42707, w42708, w42709, w42710, w42711, w42712, w42713, w42714, w42715, w42716, w42717, w42718, w42719, w42720, w42721, w42722, w42723, w42724, w42725, w42726, w42727, w42728, w42729, w42730, w42731, w42732, w42733, w42734, w42735, w42736, w42737, w42738, w42739, w42740, w42741, w42742, w42743, w42744, w42745, w42746, w42747, w42748, w42749, w42750, w42751, w42752, w42753, w42754, w42755, w42756, w42757, w42758, w42759, w42760, w42761, w42762, w42763, w42764, w42765, w42766, w42767, w42768, w42769, w42770, w42771, w42772, w42773, w42774, w42775, w42776, w42777, w42778, w42779, w42780, w42781, w42782, w42783, w42784, w42785, w42786, w42787, w42788, w42789, w42790, w42791, w42792, w42793, w42794, w42795, w42796, w42797, w42798, w42799, w42800, w42801, w42802, w42803, w42804, w42805, w42806, w42807, w42808, w42809, w42810, w42811, w42812, w42813, w42814, w42815, w42816, w42817, w42818, w42819, w42820, w42821, w42822, w42823, w42824, w42825, w42826, w42827, w42828, w42829, w42830, w42831, w42832, w42833, w42834, w42835, w42836, w42837, w42838, w42839, w42840, w42841, w42842, w42843, w42844, w42845, w42846, w42847, w42848, w42849, w42850, w42851, w42852, w42853, w42854, w42855, w42856, w42857, w42858, w42859, w42860, w42861, w42862, w42863, w42864, w42865, w42866, w42867, w42868, w42869, w42870, w42871, w42872, w42873, w42874, w42875, w42876, w42877, w42878, w42879, w42880, w42881, w42882, w42883, w42884, w42885, w42886, w42887, w42888, w42889, w42890, w42891, w42892, w42893, w42894, w42895, w42896, w42897, w42898, w42899, w42900, w42901, w42902, w42903, w42904, w42905, w42906, w42907, w42908, w42909, w42910, w42911, w42912, w42913, w42914, w42915, w42916, w42917, w42918, w42919, w42920, w42921, w42922, w42923, w42924, w42925, w42926, w42927, w42928, w42929, w42930, w42931, w42932, w42933, w42934, w42935, w42936, w42937, w42938, w42939, w42940, w42941, w42942, w42943, w42944, w42945, w42946, w42947, w42948, w42949, w42950, w42951, w42952, w42953, w42954, w42955, w42956, w42957, w42958, w42959, w42960, w42961, w42962, w42963, w42964, w42965, w42966, w42967, w42968, w42969, w42970, w42971, w42972, w42973, w42974, w42975, w42976, w42977, w42978, w42979, w42980, w42981, w42982, w42983, w42984, w42985, w42986, w42987, w42988, w42989, w42990, w42991, w42992, w42993, w42994, w42995, w42996, w42997, w42998, w42999, w43000, w43001, w43002, w43003, w43004, w43005, w43006, w43007, w43008, w43009, w43010, w43011, w43012, w43013, w43014, w43015, w43016, w43017, w43018, w43019, w43020, w43021, w43022, w43023, w43024, w43025, w43026, w43027, w43028, w43029, w43030, w43031, w43032, w43033, w43034, w43035, w43036, w43037, w43038, w43039, w43040, w43041, w43042, w43043, w43044, w43045, w43046, w43047, w43048, w43049, w43050, w43051, w43052, w43053, w43054, w43055, w43056, w43057, w43058, w43059, w43060, w43061, w43062, w43063, w43064, w43065, w43066, w43067, w43068, w43069, w43070, w43071, w43072, w43073, w43074, w43075, w43076, w43077, w43078, w43079, w43080, w43081, w43082, w43083, w43084, w43085, w43086, w43087, w43088, w43089, w43090, w43091, w43092, w43093, w43094, w43095, w43096, w43097, w43098, w43099, w43100, w43101, w43102, w43103, w43104, w43105, w43106, w43107, w43108, w43109, w43110, w43111, w43112, w43113, w43114, w43115, w43116, w43117, w43118, w43119, w43120, w43121, w43122, w43123, w43124, w43125, w43126, w43127, w43128, w43129, w43130, w43131, w43132, w43133, w43134, w43135, w43136, w43137, w43138, w43139, w43140, w43141, w43142, w43143, w43144, w43145, w43146, w43147, w43148, w43149, w43150, w43151, w43152, w43153, w43154, w43155, w43156, w43157, w43158, w43159, w43160, w43161, w43162, w43163, w43164, w43165, w43166, w43167, w43168, w43169, w43170, w43171, w43172, w43173, w43174, w43175, w43176, w43177, w43178, w43179, w43180, w43181, w43182, w43183, w43184, w43185, w43186, w43187, w43188, w43189, w43190, w43191, w43192, w43193, w43194, w43195, w43196, w43197, w43198, w43199, w43200, w43201, w43202, w43203, w43204, w43205, w43206, w43207, w43208, w43209, w43210, w43211, w43212, w43213, w43214, w43215, w43216, w43217, w43218, w43219, w43220, w43221, w43222, w43223, w43224, w43225, w43226, w43227, w43228, w43229, w43230, w43231, w43232, w43233, w43234, w43235, w43236, w43237, w43238, w43239, w43240, w43241, w43242, w43243, w43244, w43245, w43246, w43247, w43248, w43249, w43250, w43251, w43252, w43253, w43254, w43255, w43256, w43257, w43258, w43259, w43260, w43261, w43262, w43263, w43264, w43265, w43266, w43267, w43268, w43269, w43270, w43271, w43272, w43273, w43274, w43275, w43276, w43277, w43278, w43279, w43280, w43281, w43282, w43283, w43284, w43285, w43286, w43287, w43288, w43289, w43290, w43291, w43292, w43293, w43294, w43295, w43296, w43297, w43298, w43299, w43300, w43301, w43302, w43303, w43304, w43305, w43306, w43307, w43308, w43309, w43310, w43311, w43312, w43313, w43314, w43315, w43316, w43317, w43318, w43319, w43320, w43321, w43322, w43323, w43324, w43325, w43326, w43327, w43328, w43329, w43330, w43331, w43332, w43333, w43334, w43335, w43336, w43337, w43338, w43339, w43340, w43341, w43342, w43343, w43344, w43345, w43346, w43347, w43348, w43349, w43350, w43351, w43352, w43353, w43354, w43355, w43356, w43357, w43358, w43359, w43360, w43361, w43362, w43363, w43364, w43365, w43366, w43367, w43368, w43369, w43370, w43371, w43372, w43373, w43374, w43375, w43376, w43377, w43378, w43379, w43380, w43381, w43382, w43383, w43384, w43385, w43386, w43387, w43388, w43389, w43390, w43391, w43392, w43393, w43394, w43395, w43396, w43397, w43398, w43399, w43400, w43401, w43402, w43403, w43404, w43405, w43406, w43407, w43408, w43409, w43410, w43411, w43412, w43413, w43414, w43415, w43416, w43417, w43418, w43419, w43420, w43421, w43422, w43423, w43424, w43425, w43426, w43427, w43428, w43429, w43430, w43431, w43432, w43433, w43434, w43435, w43436, w43437, w43438, w43439, w43440, w43441, w43442, w43443, w43444, w43445, w43446, w43447, w43448, w43449, w43450, w43451, w43452, w43453, w43454, w43455, w43456, w43457, w43458, w43459, w43460, w43461, w43462, w43463, w43464, w43465, w43466, w43467, w43468, w43469, w43470, w43471, w43472, w43473, w43474, w43475, w43476, w43477, w43478, w43479, w43480, w43481, w43482, w43483, w43484, w43485, w43486, w43487, w43488, w43489, w43490, w43491, w43492, w43493, w43494, w43495, w43496, w43497, w43498, w43499, w43500, w43501, w43502, w43503, w43504, w43505, w43506, w43507, w43508, w43509, w43510, w43511, w43512, w43513, w43514, w43515, w43516, w43517, w43518, w43519, w43520, w43521, w43522, w43523, w43524, w43525, w43526, w43527, w43528, w43529, w43530, w43531, w43532, w43533, w43534, w43535, w43536, w43537, w43538, w43539, w43540, w43541, w43542, w43543, w43544, w43545, w43546, w43547, w43548, w43549, w43550, w43551, w43552, w43553, w43554, w43555, w43556, w43557, w43558, w43559, w43560, w43561, w43562, w43563, w43564, w43565, w43566, w43567, w43568, w43569, w43570, w43571, w43572, w43573, w43574, w43575, w43576, w43577, w43578, w43579, w43580, w43581, w43582, w43583, w43584, w43585, w43586, w43587, w43588, w43589, w43590, w43591, w43592, w43593, w43594, w43595, w43596, w43597, w43598, w43599, w43600, w43601, w43602, w43603, w43604, w43605, w43606, w43607, w43608, w43609, w43610, w43611, w43612, w43613, w43614, w43615, w43616, w43617, w43618, w43619, w43620, w43621, w43622, w43623, w43624, w43625, w43626, w43627, w43628, w43629, w43630, w43631, w43632, w43633, w43634, w43635, w43636, w43637, w43638, w43639, w43640, w43641, w43642, w43643, w43644, w43645, w43646, w43647, w43648, w43649, w43650, w43651, w43652, w43653, w43654, w43655, w43656, w43657, w43658, w43659, w43660, w43661, w43662, w43663, w43664, w43665, w43666, w43667, w43668, w43669, w43670, w43671, w43672, w43673, w43674, w43675, w43676, w43677, w43678, w43679, w43680, w43681, w43682, w43683, w43684, w43685, w43686, w43687, w43688, w43689, w43690, w43691, w43692, w43693, w43694, w43695, w43696, w43697, w43698, w43699, w43700, w43701, w43702, w43703, w43704, w43705, w43706, w43707, w43708, w43709, w43710, w43711, w43712, w43713, w43714, w43715, w43716, w43717, w43718, w43719, w43720, w43721, w43722, w43723, w43724, w43725, w43726, w43727, w43728, w43729, w43730, w43731, w43732, w43733, w43734, w43735, w43736, w43737, w43738, w43739, w43740, w43741, w43742, w43743, w43744, w43745, w43746, w43747, w43748, w43749, w43750, w43751, w43752, w43753, w43754, w43755, w43756, w43757, w43758, w43759, w43760, w43761, w43762, w43763, w43764, w43765, w43766, w43767, w43768, w43769, w43770, w43771, w43772, w43773, w43774, w43775, w43776, w43777, w43778, w43779, w43780, w43781, w43782, w43783, w43784, w43785, w43786, w43787, w43788, w43789, w43790, w43791, w43792, w43793, w43794, w43795, w43796, w43797, w43798, w43799, w43800, w43801, w43802, w43803, w43804, w43805, w43806, w43807, w43808, w43809, w43810, w43811, w43812, w43813, w43814, w43815, w43816, w43817, w43818, w43819, w43820, w43821, w43822, w43823, w43824, w43825, w43826, w43827, w43828, w43829, w43830, w43831, w43832, w43833, w43834, w43835, w43836, w43837, w43838, w43839, w43840, w43841, w43842, w43843, w43844, w43845, w43846, w43847, w43848, w43849, w43850, w43851, w43852, w43853, w43854, w43855, w43856, w43857, w43858, w43859, w43860, w43861, w43862, w43863, w43864, w43865, w43866, w43867, w43868, w43869, w43870, w43871, w43872, w43873, w43874, w43875, w43876, w43877, w43878, w43879, w43880, w43881, w43882, w43883, w43884, w43885, w43886, w43887, w43888, w43889, w43890, w43891, w43892, w43893, w43894, w43895, w43896, w43897, w43898, w43899, w43900, w43901, w43902, w43903, w43904, w43905, w43906, w43907, w43908, w43909, w43910, w43911, w43912, w43913, w43914, w43915, w43916, w43917, w43918, w43919, w43920, w43921, w43922, w43923, w43924, w43925, w43926, w43927, w43928, w43929, w43930, w43931, w43932, w43933, w43934, w43935, w43936, w43937, w43938, w43939, w43940, w43941, w43942, w43943, w43944, w43945, w43946, w43947, w43948, w43949, w43950, w43951, w43952, w43953, w43954, w43955, w43956, w43957, w43958, w43959, w43960, w43961, w43962, w43963, w43964, w43965, w43966, w43967, w43968, w43969, w43970, w43971, w43972, w43973, w43974, w43975, w43976, w43977, w43978, w43979, w43980, w43981, w43982, w43983, w43984, w43985, w43986, w43987, w43988, w43989, w43990, w43991, w43992, w43993, w43994, w43995, w43996, w43997, w43998, w43999, w44000, w44001, w44002, w44003, w44004, w44005, w44006, w44007, w44008, w44009, w44010, w44011, w44012, w44013, w44014, w44015, w44016, w44017, w44018, w44019, w44020, w44021, w44022, w44023, w44024, w44025, w44026, w44027, w44028, w44029, w44030, w44031, w44032, w44033, w44034, w44035, w44036, w44037, w44038, w44039, w44040, w44041, w44042, w44043, w44044, w44045, w44046, w44047, w44048, w44049, w44050, w44051, w44052, w44053, w44054, w44055, w44056, w44057, w44058, w44059, w44060, w44061, w44062, w44063, w44064, w44065, w44066, w44067, w44068, w44069, w44070, w44071, w44072, w44073, w44074, w44075, w44076, w44077, w44078, w44079, w44080, w44081, w44082, w44083, w44084, w44085, w44086, w44087, w44088, w44089, w44090, w44091, w44092, w44093, w44094, w44095, w44096, w44097, w44098, w44099, w44100, w44101, w44102, w44103, w44104, w44105, w44106, w44107, w44108, w44109, w44110, w44111, w44112, w44113, w44114, w44115, w44116, w44117, w44118, w44119, w44120, w44121, w44122, w44123, w44124, w44125, w44126, w44127, w44128, w44129, w44130, w44131, w44132, w44133, w44134, w44135, w44136, w44137, w44138, w44139, w44140, w44141, w44142, w44143, w44144, w44145, w44146, w44147, w44148, w44149, w44150, w44151, w44152, w44153, w44154, w44155, w44156, w44157, w44158, w44159, w44160, w44161, w44162, w44163, w44164, w44165, w44166, w44167, w44168, w44169, w44170, w44171, w44172, w44173, w44174, w44175, w44176, w44177, w44178, w44179, w44180, w44181, w44182, w44183, w44184, w44185, w44186, w44187, w44188, w44189, w44190, w44191, w44192, w44193, w44194, w44195, w44196, w44197, w44198, w44199, w44200, w44201, w44202, w44203, w44204, w44205, w44206, w44207, w44208, w44209, w44210, w44211, w44212, w44213, w44214, w44215, w44216, w44217, w44218, w44219, w44220, w44221, w44222, w44223, w44224, w44225, w44226, w44227, w44228, w44229, w44230, w44231, w44232, w44233, w44234, w44235, w44236, w44237, w44238, w44239, w44240, w44241, w44242, w44243, w44244, w44245, w44246, w44247, w44248, w44249, w44250, w44251, w44252, w44253, w44254, w44255, w44256, w44257, w44258, w44259, w44260, w44261, w44262, w44263, w44264, w44265, w44266, w44267, w44268, w44269, w44270, w44271, w44272, w44273, w44274, w44275, w44276, w44277, w44278, w44279, w44280, w44281, w44282, w44283, w44284, w44285, w44286, w44287, w44288, w44289, w44290, w44291, w44292, w44293, w44294, w44295, w44296, w44297, w44298, w44299, w44300, w44301, w44302, w44303, w44304, w44305, w44306, w44307, w44308, w44309, w44310, w44311, w44312, w44313, w44314, w44315, w44316, w44317, w44318, w44319, w44320, w44321, w44322, w44323, w44324, w44325, w44326, w44327, w44328, w44329, w44330, w44331, w44332, w44333, w44334, w44335, w44336, w44337, w44338, w44339, w44340, w44341, w44342, w44343, w44344, w44345, w44346, w44347, w44348, w44349, w44350, w44351, w44352, w44353, w44354, w44355, w44356, w44357, w44358, w44359, w44360, w44361, w44362, w44363, w44364, w44365, w44366, w44367, w44368, w44369, w44370, w44371, w44372, w44373, w44374, w44375, w44376, w44377, w44378, w44379, w44380, w44381, w44382, w44383, w44384, w44385, w44386, w44387, w44388, w44389, w44390, w44391, w44392, w44393, w44394, w44395, w44396, w44397, w44398, w44399, w44400, w44401, w44402, w44403, w44404, w44405, w44406, w44407, w44408, w44409, w44410, w44411, w44412, w44413, w44414, w44415, w44416, w44417, w44418, w44419, w44420, w44421, w44422, w44423, w44424, w44425, w44426, w44427, w44428, w44429, w44430, w44431, w44432, w44433, w44434, w44435, w44436, w44437, w44438, w44439, w44440, w44441, w44442, w44443, w44444, w44445, w44446, w44447, w44448, w44449, w44450, w44451, w44452, w44453, w44454, w44455, w44456, w44457, w44458, w44459, w44460, w44461, w44462, w44463, w44464, w44465, w44466, w44467, w44468, w44469, w44470, w44471, w44472, w44473, w44474, w44475, w44476, w44477, w44478, w44479, w44480, w44481, w44482, w44483, w44484, w44485, w44486, w44487, w44488, w44489, w44490, w44491, w44492, w44493, w44494, w44495, w44496, w44497, w44498, w44499, w44500, w44501, w44502, w44503, w44504, w44505, w44506, w44507, w44508, w44509, w44510, w44511, w44512, w44513, w44514, w44515, w44516, w44517, w44518, w44519, w44520, w44521, w44522, w44523, w44524, w44525, w44526, w44527, w44528, w44529, w44530, w44531, w44532, w44533, w44534, w44535, w44536, w44537, w44538, w44539, w44540, w44541, w44542, w44543, w44544, w44545, w44546, w44547, w44548, w44549, w44550, w44551, w44552, w44553, w44554, w44555, w44556, w44557, w44558, w44559, w44560, w44561, w44562, w44563, w44564, w44565, w44566, w44567, w44568, w44569, w44570, w44571, w44572, w44573, w44574, w44575, w44576, w44577, w44578, w44579, w44580, w44581, w44582, w44583, w44584, w44585, w44586, w44587, w44588, w44589, w44590, w44591, w44592, w44593, w44594, w44595, w44596, w44597, w44598, w44599, w44600, w44601, w44602, w44603, w44604, w44605, w44606, w44607, w44608, w44609, w44610, w44611, w44612, w44613, w44614, w44615, w44616, w44617, w44618, w44619, w44620, w44621, w44622, w44623, w44624, w44625, w44626, w44627, w44628, w44629, w44630, w44631, w44632, w44633, w44634, w44635, w44636, w44637, w44638, w44639, w44640, w44641, w44642, w44643, w44644, w44645, w44646, w44647, w44648, w44649, w44650, w44651, w44652, w44653, w44654, w44655, w44656, w44657, w44658, w44659, w44660, w44661, w44662, w44663, w44664, w44665, w44666, w44667, w44668, w44669, w44670, w44671, w44672, w44673, w44674, w44675, w44676, w44677, w44678, w44679, w44680, w44681, w44682, w44683, w44684, w44685, w44686, w44687, w44688, w44689, w44690, w44691, w44692, w44693, w44694, w44695, w44696, w44697, w44698, w44699, w44700, w44701, w44702, w44703, w44704, w44705, w44706, w44707, w44708, w44709, w44710, w44711, w44712, w44713, w44714, w44715, w44716, w44717, w44718, w44719, w44720, w44721, w44722, w44723, w44724, w44725, w44726, w44727, w44728, w44729, w44730, w44731, w44732, w44733, w44734, w44735, w44736, w44737, w44738, w44739, w44740, w44741, w44742, w44743, w44744, w44745, w44746, w44747, w44748, w44749, w44750, w44751, w44752, w44753, w44754, w44755, w44756, w44757, w44758, w44759, w44760, w44761, w44762, w44763, w44764, w44765, w44766, w44767, w44768, w44769, w44770, w44771, w44772, w44773, w44774, w44775, w44776, w44777, w44778, w44779, w44780, w44781, w44782, w44783, w44784, w44785, w44786, w44787, w44788, w44789, w44790, w44791, w44792, w44793, w44794, w44795, w44796, w44797, w44798, w44799, w44800, w44801, w44802, w44803, w44804, w44805, w44806, w44807, w44808, w44809, w44810, w44811, w44812, w44813, w44814, w44815, w44816, w44817, w44818, w44819, w44820, w44821, w44822, w44823, w44824, w44825, w44826, w44827, w44828, w44829, w44830, w44831, w44832, w44833, w44834, w44835, w44836, w44837, w44838, w44839, w44840, w44841, w44842, w44843, w44844, w44845, w44846, w44847, w44848, w44849, w44850, w44851, w44852, w44853, w44854, w44855, w44856, w44857, w44858, w44859, w44860, w44861, w44862, w44863, w44864, w44865, w44866, w44867, w44868, w44869, w44870, w44871, w44872, w44873, w44874, w44875, w44876, w44877, w44878, w44879, w44880, w44881, w44882, w44883, w44884, w44885, w44886, w44887, w44888, w44889, w44890, w44891, w44892, w44893, w44894, w44895, w44896, w44897, w44898, w44899, w44900, w44901, w44902, w44903, w44904, w44905, w44906, w44907, w44908, w44909, w44910, w44911, w44912, w44913, w44914, w44915, w44916, w44917, w44918, w44919, w44920, w44921, w44922, w44923, w44924, w44925, w44926, w44927, w44928, w44929, w44930, w44931, w44932, w44933, w44934, w44935, w44936, w44937, w44938, w44939, w44940, w44941, w44942, w44943, w44944, w44945, w44946, w44947, w44948, w44949, w44950, w44951, w44952, w44953, w44954, w44955, w44956, w44957, w44958, w44959, w44960, w44961, w44962, w44963, w44964, w44965, w44966, w44967, w44968, w44969, w44970, w44971, w44972, w44973, w44974, w44975, w44976, w44977, w44978, w44979, w44980, w44981, w44982, w44983, w44984, w44985, w44986, w44987, w44988, w44989, w44990, w44991, w44992, w44993, w44994, w44995, w44996, w44997, w44998, w44999, w45000, w45001, w45002, w45003, w45004, w45005, w45006, w45007, w45008, w45009, w45010, w45011, w45012, w45013, w45014, w45015, w45016, w45017, w45018, w45019, w45020, w45021, w45022, w45023, w45024, w45025, w45026, w45027, w45028, w45029, w45030, w45031, w45032, w45033, w45034, w45035, w45036, w45037, w45038, w45039, w45040, w45041, w45042, w45043, w45044, w45045, w45046, w45047, w45048, w45049, w45050, w45051, w45052, w45053, w45054, w45055, w45056, w45057, w45058, w45059, w45060, w45061, w45062, w45063, w45064, w45065, w45066, w45067, w45068, w45069, w45070, w45071, w45072, w45073, w45074, w45075, w45076, w45077, w45078, w45079, w45080, w45081, w45082, w45083, w45084, w45085, w45086, w45087, w45088, w45089, w45090, w45091, w45092, w45093, w45094, w45095, w45096, w45097, w45098, w45099, w45100, w45101, w45102, w45103, w45104, w45105, w45106, w45107, w45108, w45109, w45110, w45111, w45112, w45113, w45114, w45115, w45116, w45117, w45118, w45119, w45120, w45121, w45122, w45123, w45124, w45125, w45126, w45127, w45128, w45129, w45130, w45131, w45132, w45133, w45134, w45135, w45136, w45137, w45138, w45139, w45140, w45141, w45142, w45143, w45144, w45145, w45146, w45147, w45148, w45149, w45150, w45151, w45152, w45153, w45154, w45155, w45156, w45157, w45158, w45159, w45160, w45161, w45162, w45163, w45164, w45165, w45166, w45167, w45168, w45169, w45170, w45171, w45172, w45173, w45174, w45175, w45176, w45177, w45178, w45179, w45180, w45181, w45182, w45183, w45184, w45185, w45186, w45187, w45188, w45189, w45190, w45191, w45192, w45193, w45194, w45195, w45196, w45197, w45198, w45199, w45200, w45201, w45202, w45203, w45204, w45205, w45206, w45207, w45208, w45209, w45210, w45211, w45212, w45213, w45214, w45215, w45216, w45217, w45218, w45219, w45220, w45221, w45222, w45223, w45224, w45225, w45226, w45227, w45228, w45229, w45230, w45231, w45232, w45233, w45234, w45235, w45236, w45237, w45238, w45239, w45240, w45241, w45242, w45243, w45244, w45245, w45246, w45247, w45248, w45249, w45250, w45251, w45252, w45253, w45254, w45255, w45256, w45257, w45258, w45259, w45260, w45261, w45262, w45263, w45264, w45265, w45266, w45267, w45268, w45269, w45270, w45271, w45272, w45273, w45274, w45275, w45276, w45277, w45278, w45279, w45280, w45281, w45282, w45283, w45284, w45285, w45286, w45287, w45288, w45289, w45290, w45291, w45292, w45293, w45294, w45295, w45296, w45297, w45298, w45299, w45300, w45301, w45302, w45303, w45304, w45305, w45306, w45307, w45308, w45309, w45310, w45311, w45312, w45313, w45314, w45315, w45316, w45317, w45318, w45319, w45320, w45321, w45322, w45323, w45324, w45325, w45326, w45327, w45328, w45329, w45330, w45331, w45332, w45333, w45334, w45335, w45336, w45337, w45338, w45339, w45340, w45341, w45342, w45343, w45344, w45345, w45346, w45347, w45348, w45349, w45350, w45351, w45352, w45353, w45354, w45355, w45356, w45357, w45358, w45359, w45360, w45361, w45362, w45363, w45364, w45365, w45366, w45367, w45368, w45369, w45370, w45371, w45372, w45373, w45374, w45375, w45376, w45377, w45378, w45379, w45380, w45381, w45382, w45383, w45384, w45385, w45386, w45387, w45388, w45389, w45390, w45391, w45392, w45393, w45394, w45395, w45396, w45397, w45398, w45399, w45400, w45401, w45402, w45403, w45404, w45405, w45406, w45407, w45408, w45409, w45410, w45411, w45412, w45413, w45414, w45415, w45416, w45417, w45418, w45419, w45420, w45421, w45422, w45423, w45424, w45425, w45426, w45427, w45428, w45429, w45430, w45431, w45432, w45433, w45434, w45435, w45436, w45437, w45438, w45439, w45440, w45441, w45442, w45443, w45444, w45445, w45446, w45447, w45448, w45449, w45450, w45451, w45452, w45453, w45454, w45455, w45456, w45457, w45458, w45459, w45460, w45461, w45462, w45463, w45464, w45465, w45466, w45467, w45468, w45469, w45470, w45471, w45472, w45473, w45474, w45475, w45476, w45477, w45478, w45479, w45480, w45481, w45482, w45483, w45484, w45485, w45486, w45487, w45488, w45489, w45490, w45491, w45492, w45493, w45494, w45495, w45496, w45497, w45498, w45499, w45500, w45501, w45502, w45503, w45504, w45505, w45506, w45507, w45508, w45509, w45510, w45511, w45512, w45513, w45514, w45515, w45516, w45517, w45518, w45519, w45520, w45521, w45522, w45523, w45524, w45525, w45526, w45527, w45528, w45529, w45530, w45531, w45532, w45533, w45534, w45535, w45536, w45537, w45538, w45539, w45540, w45541, w45542, w45543, w45544, w45545, w45546, w45547, w45548, w45549, w45550, w45551, w45552, w45553, w45554, w45555, w45556, w45557, w45558, w45559, w45560, w45561, w45562, w45563, w45564, w45565, w45566, w45567, w45568, w45569, w45570, w45571, w45572, w45573, w45574, w45575, w45576, w45577, w45578, w45579, w45580, w45581, w45582, w45583, w45584, w45585, w45586, w45587, w45588, w45589, w45590, w45591, w45592, w45593, w45594, w45595, w45596, w45597, w45598, w45599, w45600, w45601, w45602, w45603, w45604, w45605, w45606, w45607, w45608, w45609, w45610, w45611, w45612, w45613, w45614, w45615, w45616, w45617, w45618, w45619, w45620, w45621, w45622, w45623, w45624, w45625, w45626, w45627, w45628, w45629, w45630, w45631, w45632, w45633, w45634, w45635, w45636, w45637, w45638, w45639, w45640, w45641, w45642, w45643, w45644, w45645, w45646, w45647, w45648, w45649, w45650, w45651, w45652, w45653, w45654, w45655, w45656, w45657, w45658, w45659, w45660, w45661, w45662, w45663, w45664, w45665, w45666, w45667, w45668, w45669, w45670, w45671, w45672, w45673, w45674, w45675, w45676, w45677, w45678, w45679, w45680, w45681, w45682, w45683, w45684, w45685, w45686, w45687, w45688, w45689, w45690, w45691, w45692, w45693, w45694, w45695, w45696, w45697, w45698, w45699, w45700, w45701, w45702, w45703, w45704, w45705, w45706, w45707, w45708, w45709, w45710, w45711, w45712, w45713, w45714, w45715, w45716, w45717, w45718, w45719, w45720, w45721, w45722, w45723, w45724, w45725, w45726, w45727, w45728, w45729, w45730, w45731, w45732, w45733, w45734, w45735, w45736, w45737, w45738, w45739, w45740, w45741, w45742, w45743, w45744, w45745, w45746, w45747, w45748, w45749, w45750, w45751, w45752, w45753, w45754, w45755, w45756, w45757, w45758, w45759, w45760, w45761, w45762, w45763, w45764, w45765, w45766, w45767, w45768, w45769, w45770, w45771, w45772, w45773, w45774, w45775, w45776, w45777, w45778, w45779, w45780, w45781, w45782, w45783, w45784, w45785, w45786, w45787, w45788, w45789, w45790, w45791, w45792, w45793, w45794, w45795, w45796, w45797, w45798, w45799, w45800, w45801, w45802, w45803, w45804, w45805, w45806, w45807, w45808, w45809, w45810, w45811, w45812, w45813, w45814, w45815, w45816, w45817, w45818, w45819, w45820, w45821, w45822, w45823, w45824, w45825, w45826, w45827, w45828, w45829, w45830, w45831, w45832, w45833, w45834, w45835, w45836, w45837, w45838, w45839, w45840, w45841, w45842, w45843, w45844, w45845, w45846, w45847, w45848, w45849, w45850, w45851, w45852, w45853, w45854, w45855, w45856, w45857, w45858, w45859, w45860, w45861, w45862, w45863, w45864, w45865, w45866, w45867, w45868, w45869, w45870, w45871, w45872, w45873, w45874, w45875, w45876, w45877, w45878, w45879, w45880, w45881, w45882, w45883, w45884, w45885, w45886, w45887, w45888, w45889, w45890, w45891, w45892, w45893, w45894, w45895, w45896, w45897, w45898, w45899, w45900, w45901, w45902, w45903, w45904, w45905, w45906, w45907, w45908, w45909, w45910, w45911, w45912, w45913, w45914, w45915, w45916, w45917, w45918, w45919, w45920, w45921, w45922, w45923, w45924, w45925, w45926, w45927, w45928, w45929, w45930, w45931, w45932, w45933, w45934, w45935, w45936, w45937, w45938, w45939, w45940, w45941, w45942, w45943, w45944, w45945, w45946, w45947, w45948, w45949, w45950, w45951, w45952, w45953, w45954, w45955, w45956, w45957, w45958, w45959, w45960, w45961, w45962, w45963, w45964, w45965, w45966, w45967, w45968, w45969, w45970, w45971, w45972, w45973, w45974, w45975, w45976, w45977, w45978, w45979, w45980, w45981, w45982, w45983, w45984, w45985, w45986, w45987, w45988, w45989, w45990, w45991, w45992, w45993, w45994, w45995, w45996, w45997, w45998, w45999, w46000, w46001, w46002, w46003, w46004, w46005, w46006, w46007, w46008, w46009, w46010, w46011, w46012, w46013, w46014, w46015, w46016, w46017, w46018, w46019, w46020, w46021, w46022, w46023, w46024, w46025, w46026, w46027, w46028, w46029, w46030, w46031, w46032, w46033, w46034, w46035, w46036, w46037, w46038, w46039, w46040, w46041, w46042, w46043, w46044, w46045, w46046, w46047, w46048, w46049, w46050, w46051, w46052, w46053, w46054, w46055, w46056, w46057, w46058, w46059, w46060, w46061, w46062, w46063, w46064, w46065, w46066, w46067, w46068, w46069, w46070, w46071, w46072, w46073, w46074, w46075, w46076, w46077, w46078, w46079, w46080, w46081, w46082, w46083, w46084, w46085, w46086, w46087, w46088, w46089, w46090, w46091, w46092, w46093, w46094, w46095, w46096, w46097, w46098, w46099, w46100, w46101, w46102, w46103, w46104, w46105, w46106, w46107, w46108, w46109, w46110, w46111, w46112, w46113, w46114, w46115, w46116, w46117, w46118, w46119, w46120, w46121, w46122, w46123, w46124, w46125, w46126, w46127, w46128, w46129, w46130, w46131, w46132, w46133, w46134, w46135, w46136, w46137, w46138, w46139, w46140, w46141, w46142, w46143, w46144, w46145, w46146, w46147, w46148, w46149, w46150, w46151, w46152, w46153, w46154, w46155, w46156, w46157, w46158, w46159, w46160, w46161, w46162, w46163, w46164, w46165, w46166, w46167, w46168, w46169, w46170, w46171, w46172, w46173, w46174, w46175, w46176, w46177, w46178, w46179, w46180, w46181, w46182, w46183, w46184, w46185, w46186, w46187, w46188, w46189, w46190, w46191, w46192, w46193, w46194, w46195, w46196, w46197, w46198, w46199, w46200, w46201, w46202, w46203, w46204, w46205, w46206, w46207, w46208, w46209, w46210, w46211, w46212, w46213, w46214, w46215, w46216, w46217, w46218, w46219, w46220, w46221, w46222, w46223, w46224, w46225, w46226, w46227, w46228, w46229, w46230, w46231, w46232, w46233, w46234, w46235, w46236, w46237, w46238, w46239, w46240, w46241, w46242, w46243, w46244, w46245, w46246, w46247, w46248, w46249, w46250, w46251, w46252, w46253, w46254, w46255, w46256, w46257, w46258, w46259, w46260, w46261, w46262, w46263, w46264, w46265, w46266, w46267, w46268, w46269, w46270, w46271, w46272, w46273, w46274, w46275, w46276, w46277, w46278, w46279, w46280, w46281, w46282, w46283, w46284, w46285, w46286, w46287, w46288, w46289, w46290, w46291, w46292, w46293, w46294, w46295, w46296, w46297, w46298, w46299, w46300, w46301, w46302, w46303, w46304, w46305, w46306, w46307, w46308, w46309, w46310, w46311, w46312, w46313, w46314, w46315, w46316, w46317, w46318, w46319, w46320, w46321, w46322, w46323, w46324, w46325, w46326, w46327, w46328, w46329, w46330, w46331, w46332, w46333, w46334, w46335, w46336, w46337, w46338, w46339, w46340, w46341, w46342, w46343, w46344, w46345, w46346, w46347, w46348, w46349, w46350, w46351, w46352, w46353, w46354, w46355, w46356, w46357, w46358, w46359, w46360, w46361, w46362, w46363, w46364, w46365, w46366, w46367, w46368, w46369, w46370, w46371, w46372, w46373, w46374, w46375, w46376, w46377, w46378, w46379, w46380, w46381, w46382, w46383, w46384, w46385, w46386, w46387, w46388, w46389, w46390, w46391, w46392, w46393, w46394, w46395, w46396, w46397, w46398, w46399, w46400, w46401, w46402, w46403, w46404, w46405, w46406, w46407, w46408, w46409, w46410, w46411, w46412, w46413, w46414, w46415, w46416, w46417, w46418, w46419, w46420, w46421, w46422, w46423, w46424, w46425, w46426, w46427, w46428, w46429, w46430, w46431, w46432, w46433, w46434, w46435, w46436, w46437, w46438, w46439, w46440, w46441, w46442, w46443, w46444, w46445, w46446, w46447, w46448, w46449, w46450, w46451, w46452, w46453, w46454, w46455, w46456, w46457, w46458, w46459, w46460, w46461, w46462, w46463, w46464, w46465, w46466, w46467, w46468, w46469, w46470, w46471, w46472, w46473, w46474, w46475, w46476, w46477, w46478, w46479, w46480, w46481, w46482, w46483, w46484, w46485, w46486, w46487, w46488, w46489, w46490, w46491, w46492, w46493, w46494, w46495, w46496, w46497, w46498, w46499, w46500, w46501, w46502, w46503, w46504, w46505, w46506, w46507, w46508, w46509, w46510, w46511, w46512, w46513, w46514, w46515, w46516, w46517, w46518, w46519, w46520, w46521, w46522, w46523, w46524, w46525, w46526, w46527, w46528, w46529, w46530, w46531, w46532, w46533, w46534, w46535, w46536, w46537, w46538, w46539, w46540, w46541, w46542, w46543, w46544, w46545, w46546, w46547, w46548, w46549, w46550, w46551, w46552, w46553, w46554, w46555, w46556, w46557, w46558, w46559, w46560, w46561, w46562, w46563, w46564, w46565, w46566, w46567, w46568, w46569, w46570, w46571, w46572, w46573, w46574, w46575, w46576, w46577, w46578, w46579, w46580, w46581, w46582, w46583, w46584, w46585, w46586, w46587, w46588, w46589, w46590, w46591, w46592, w46593, w46594, w46595, w46596, w46597, w46598, w46599, w46600, w46601, w46602, w46603, w46604, w46605, w46606, w46607, w46608, w46609, w46610, w46611, w46612, w46613, w46614, w46615, w46616, w46617, w46618, w46619, w46620, w46621, w46622, w46623, w46624, w46625, w46626, w46627, w46628, w46629, w46630, w46631, w46632, w46633, w46634, w46635, w46636, w46637, w46638, w46639, w46640, w46641, w46642, w46643, w46644, w46645, w46646, w46647, w46648, w46649, w46650, w46651, w46652, w46653, w46654, w46655, w46656, w46657, w46658, w46659, w46660, w46661, w46662, w46663, w46664, w46665, w46666, w46667, w46668, w46669, w46670, w46671, w46672, w46673, w46674, w46675, w46676, w46677, w46678, w46679, w46680, w46681, w46682, w46683, w46684, w46685, w46686, w46687, w46688, w46689, w46690, w46691, w46692, w46693, w46694, w46695, w46696, w46697, w46698, w46699, w46700, w46701, w46702, w46703, w46704, w46705, w46706, w46707, w46708, w46709, w46710, w46711, w46712, w46713, w46714, w46715, w46716, w46717, w46718, w46719, w46720, w46721, w46722, w46723, w46724, w46725, w46726, w46727, w46728, w46729, w46730, w46731, w46732, w46733, w46734, w46735, w46736, w46737, w46738, w46739, w46740, w46741, w46742, w46743, w46744, w46745, w46746, w46747, w46748, w46749, w46750, w46751, w46752, w46753, w46754, w46755, w46756, w46757, w46758, w46759, w46760, w46761, w46762, w46763, w46764, w46765, w46766, w46767, w46768, w46769, w46770, w46771, w46772, w46773, w46774, w46775, w46776, w46777, w46778, w46779, w46780, w46781, w46782, w46783, w46784, w46785, w46786, w46787, w46788, w46789, w46790, w46791, w46792, w46793, w46794, w46795, w46796, w46797, w46798, w46799, w46800, w46801, w46802, w46803, w46804, w46805, w46806, w46807, w46808, w46809, w46810, w46811, w46812, w46813, w46814, w46815, w46816, w46817, w46818, w46819, w46820, w46821, w46822, w46823, w46824, w46825, w46826, w46827, w46828, w46829, w46830, w46831, w46832, w46833, w46834, w46835, w46836, w46837, w46838, w46839, w46840, w46841, w46842, w46843, w46844, w46845, w46846, w46847, w46848, w46849, w46850, w46851, w46852, w46853, w46854, w46855, w46856, w46857, w46858, w46859, w46860, w46861, w46862, w46863, w46864, w46865, w46866, w46867, w46868, w46869, w46870, w46871, w46872, w46873, w46874, w46875, w46876, w46877, w46878, w46879, w46880, w46881, w46882, w46883, w46884, w46885, w46886, w46887, w46888, w46889, w46890, w46891, w46892, w46893, w46894, w46895, w46896, w46897, w46898, w46899, w46900, w46901, w46902, w46903, w46904, w46905, w46906, w46907, w46908, w46909, w46910, w46911, w46912, w46913, w46914, w46915, w46916, w46917, w46918, w46919, w46920, w46921, w46922, w46923, w46924, w46925, w46926, w46927, w46928, w46929, w46930, w46931, w46932, w46933, w46934, w46935, w46936, w46937, w46938, w46939, w46940, w46941, w46942, w46943, w46944, w46945, w46946, w46947, w46948, w46949, w46950, w46951, w46952, w46953, w46954, w46955, w46956, w46957, w46958, w46959, w46960, w46961, w46962, w46963, w46964, w46965, w46966, w46967, w46968, w46969, w46970, w46971, w46972, w46973, w46974, w46975, w46976, w46977, w46978, w46979, w46980, w46981, w46982, w46983, w46984, w46985, w46986, w46987, w46988, w46989, w46990, w46991, w46992, w46993, w46994, w46995, w46996, w46997, w46998, w46999, w47000, w47001, w47002, w47003, w47004, w47005, w47006, w47007, w47008, w47009, w47010, w47011, w47012, w47013, w47014, w47015, w47016, w47017, w47018, w47019, w47020, w47021, w47022, w47023, w47024, w47025, w47026, w47027, w47028, w47029, w47030, w47031, w47032, w47033, w47034, w47035, w47036, w47037, w47038, w47039, w47040, w47041, w47042, w47043, w47044, w47045, w47046, w47047, w47048, w47049, w47050, w47051, w47052, w47053, w47054, w47055, w47056, w47057, w47058, w47059, w47060, w47061, w47062, w47063, w47064, w47065, w47066, w47067, w47068, w47069, w47070, w47071, w47072, w47073, w47074, w47075, w47076, w47077, w47078, w47079, w47080, w47081, w47082, w47083, w47084, w47085, w47086, w47087, w47088, w47089, w47090, w47091, w47092, w47093, w47094, w47095, w47096, w47097, w47098, w47099, w47100, w47101, w47102, w47103, w47104, w47105, w47106, w47107, w47108, w47109, w47110, w47111, w47112, w47113, w47114, w47115, w47116, w47117, w47118, w47119, w47120, w47121, w47122, w47123, w47124, w47125, w47126, w47127, w47128, w47129, w47130, w47131, w47132, w47133, w47134, w47135, w47136, w47137, w47138, w47139, w47140, w47141, w47142, w47143, w47144, w47145, w47146, w47147, w47148, w47149, w47150, w47151, w47152, w47153, w47154, w47155, w47156, w47157, w47158, w47159, w47160, w47161, w47162, w47163, w47164, w47165, w47166, w47167, w47168, w47169, w47170, w47171, w47172, w47173, w47174, w47175, w47176, w47177, w47178, w47179, w47180, w47181, w47182, w47183, w47184, w47185, w47186, w47187, w47188, w47189, w47190, w47191, w47192, w47193, w47194, w47195, w47196, w47197, w47198, w47199, w47200, w47201, w47202, w47203, w47204, w47205, w47206, w47207, w47208, w47209, w47210, w47211, w47212, w47213, w47214, w47215, w47216, w47217, w47218, w47219, w47220, w47221, w47222, w47223, w47224, w47225, w47226, w47227, w47228, w47229, w47230, w47231, w47232, w47233, w47234, w47235, w47236, w47237, w47238, w47239, w47240, w47241, w47242, w47243, w47244, w47245, w47246, w47247, w47248, w47249, w47250, w47251, w47252, w47253, w47254, w47255, w47256, w47257, w47258, w47259, w47260, w47261, w47262, w47263, w47264, w47265, w47266, w47267, w47268, w47269, w47270, w47271, w47272, w47273, w47274, w47275, w47276, w47277, w47278, w47279, w47280, w47281, w47282, w47283, w47284, w47285, w47286, w47287, w47288, w47289, w47290, w47291, w47292, w47293, w47294, w47295, w47296, w47297, w47298, w47299, w47300, w47301, w47302, w47303, w47304, w47305, w47306, w47307, w47308, w47309, w47310, w47311, w47312, w47313, w47314, w47315, w47316, w47317, w47318, w47319, w47320, w47321, w47322, w47323, w47324, w47325, w47326, w47327, w47328, w47329, w47330, w47331, w47332, w47333, w47334, w47335, w47336, w47337, w47338, w47339, w47340, w47341, w47342, w47343, w47344, w47345, w47346, w47347, w47348, w47349, w47350, w47351, w47352, w47353, w47354, w47355, w47356, w47357, w47358, w47359, w47360, w47361, w47362, w47363, w47364, w47365, w47366, w47367, w47368, w47369, w47370, w47371, w47372, w47373, w47374, w47375, w47376, w47377, w47378, w47379, w47380, w47381, w47382, w47383, w47384, w47385, w47386, w47387, w47388, w47389, w47390, w47391, w47392, w47393, w47394, w47395, w47396, w47397, w47398, w47399, w47400, w47401, w47402, w47403, w47404, w47405, w47406, w47407, w47408, w47409, w47410, w47411, w47412, w47413, w47414, w47415, w47416, w47417, w47418, w47419, w47420, w47421, w47422, w47423, w47424, w47425, w47426, w47427, w47428, w47429, w47430, w47431, w47432, w47433, w47434, w47435, w47436, w47437, w47438, w47439, w47440, w47441, w47442, w47443, w47444, w47445, w47446, w47447, w47448, w47449, w47450, w47451, w47452, w47453, w47454, w47455, w47456, w47457, w47458, w47459, w47460, w47461, w47462, w47463, w47464, w47465, w47466, w47467, w47468, w47469, w47470, w47471, w47472, w47473, w47474, w47475, w47476, w47477, w47478, w47479, w47480, w47481, w47482, w47483, w47484, w47485, w47486, w47487, w47488, w47489, w47490, w47491, w47492, w47493, w47494, w47495, w47496, w47497, w47498, w47499, w47500, w47501, w47502, w47503, w47504, w47505, w47506, w47507, w47508, w47509, w47510, w47511, w47512, w47513, w47514, w47515, w47516, w47517, w47518, w47519, w47520, w47521, w47522, w47523, w47524, w47525, w47526, w47527, w47528, w47529, w47530, w47531, w47532, w47533, w47534, w47535, w47536, w47537, w47538, w47539, w47540, w47541, w47542, w47543, w47544, w47545, w47546, w47547, w47548, w47549, w47550, w47551, w47552, w47553, w47554, w47555, w47556, w47557, w47558, w47559, w47560, w47561, w47562, w47563, w47564, w47565, w47566, w47567, w47568, w47569, w47570, w47571, w47572, w47573, w47574, w47575, w47576, w47577, w47578, w47579, w47580, w47581, w47582, w47583, w47584, w47585, w47586, w47587, w47588, w47589, w47590, w47591, w47592, w47593, w47594, w47595, w47596, w47597, w47598, w47599, w47600, w47601, w47602, w47603, w47604, w47605, w47606, w47607, w47608, w47609, w47610, w47611, w47612, w47613, w47614, w47615, w47616, w47617, w47618, w47619, w47620, w47621, w47622, w47623, w47624, w47625, w47626, w47627, w47628, w47629, w47630, w47631, w47632, w47633, w47634, w47635, w47636, w47637, w47638, w47639, w47640, w47641, w47642, w47643, w47644, w47645, w47646, w47647, w47648, w47649, w47650, w47651, w47652, w47653, w47654, w47655, w47656, w47657, w47658, w47659, w47660, w47661, w47662, w47663, w47664, w47665, w47666, w47667, w47668, w47669, w47670, w47671, w47672, w47673, w47674, w47675, w47676, w47677, w47678, w47679, w47680, w47681, w47682, w47683, w47684, w47685, w47686, w47687, w47688, w47689, w47690, w47691, w47692, w47693, w47694, w47695, w47696, w47697, w47698, w47699, w47700, w47701, w47702, w47703, w47704, w47705, w47706, w47707, w47708, w47709, w47710, w47711, w47712, w47713, w47714, w47715, w47716, w47717, w47718, w47719, w47720, w47721, w47722, w47723, w47724, w47725, w47726, w47727, w47728, w47729, w47730, w47731, w47732, w47733, w47734, w47735, w47736, w47737, w47738, w47739, w47740, w47741, w47742, w47743, w47744, w47745, w47746, w47747, w47748, w47749, w47750, w47751, w47752, w47753, w47754, w47755, w47756, w47757, w47758, w47759, w47760, w47761, w47762, w47763, w47764, w47765, w47766, w47767, w47768, w47769, w47770, w47771, w47772, w47773, w47774, w47775, w47776, w47777, w47778, w47779, w47780, w47781, w47782, w47783, w47784, w47785, w47786, w47787, w47788, w47789, w47790, w47791, w47792, w47793, w47794, w47795, w47796, w47797, w47798, w47799, w47800, w47801, w47802, w47803, w47804, w47805, w47806, w47807, w47808, w47809, w47810, w47811, w47812, w47813, w47814, w47815, w47816, w47817, w47818, w47819, w47820, w47821, w47822, w47823, w47824, w47825, w47826, w47827, w47828, w47829, w47830, w47831, w47832, w47833, w47834, w47835, w47836, w47837, w47838, w47839, w47840, w47841, w47842, w47843, w47844, w47845, w47846, w47847, w47848, w47849, w47850, w47851, w47852, w47853, w47854, w47855, w47856, w47857, w47858, w47859, w47860, w47861, w47862, w47863, w47864, w47865, w47866, w47867, w47868, w47869, w47870, w47871, w47872, w47873, w47874, w47875, w47876, w47877, w47878, w47879, w47880, w47881, w47882, w47883, w47884, w47885, w47886, w47887, w47888, w47889, w47890, w47891, w47892, w47893, w47894, w47895, w47896, w47897, w47898, w47899, w47900, w47901, w47902, w47903, w47904, w47905, w47906, w47907, w47908, w47909, w47910, w47911, w47912, w47913, w47914, w47915, w47916, w47917, w47918, w47919, w47920, w47921, w47922, w47923, w47924, w47925, w47926, w47927, w47928, w47929, w47930, w47931, w47932, w47933, w47934, w47935, w47936, w47937, w47938, w47939, w47940, w47941, w47942, w47943, w47944, w47945, w47946, w47947, w47948, w47949, w47950, w47951, w47952, w47953, w47954, w47955, w47956, w47957, w47958, w47959, w47960, w47961, w47962, w47963, w47964, w47965, w47966, w47967, w47968, w47969, w47970, w47971, w47972, w47973, w47974, w47975, w47976, w47977, w47978, w47979, w47980, w47981, w47982, w47983, w47984, w47985, w47986, w47987, w47988, w47989, w47990, w47991, w47992, w47993, w47994, w47995, w47996, w47997, w47998, w47999, w48000, w48001, w48002, w48003, w48004, w48005, w48006, w48007, w48008, w48009, w48010, w48011, w48012, w48013, w48014, w48015, w48016, w48017, w48018, w48019, w48020, w48021, w48022, w48023, w48024, w48025, w48026, w48027, w48028, w48029, w48030, w48031, w48032, w48033, w48034, w48035, w48036, w48037, w48038, w48039, w48040, w48041, w48042, w48043, w48044, w48045, w48046, w48047, w48048, w48049, w48050, w48051, w48052, w48053, w48054, w48055, w48056, w48057, w48058, w48059, w48060, w48061, w48062, w48063, w48064, w48065, w48066, w48067, w48068, w48069, w48070, w48071, w48072, w48073, w48074, w48075, w48076, w48077, w48078, w48079, w48080, w48081, w48082, w48083, w48084, w48085, w48086, w48087, w48088, w48089, w48090, w48091, w48092, w48093, w48094, w48095, w48096, w48097, w48098, w48099, w48100, w48101, w48102, w48103, w48104, w48105, w48106, w48107, w48108, w48109, w48110, w48111, w48112, w48113, w48114, w48115, w48116, w48117, w48118, w48119, w48120, w48121, w48122, w48123, w48124, w48125, w48126, w48127, w48128, w48129, w48130, w48131, w48132, w48133, w48134, w48135, w48136, w48137, w48138, w48139, w48140, w48141, w48142, w48143, w48144, w48145, w48146, w48147, w48148, w48149, w48150, w48151, w48152, w48153, w48154, w48155, w48156, w48157, w48158, w48159, w48160, w48161, w48162, w48163, w48164, w48165, w48166, w48167, w48168, w48169, w48170, w48171, w48172, w48173, w48174, w48175, w48176, w48177, w48178, w48179, w48180, w48181, w48182, w48183, w48184, w48185, w48186, w48187, w48188, w48189, w48190, w48191, w48192, w48193, w48194, w48195, w48196, w48197, w48198, w48199, w48200, w48201, w48202, w48203, w48204, w48205, w48206, w48207, w48208, w48209, w48210, w48211, w48212, w48213, w48214, w48215, w48216, w48217, w48218, w48219, w48220, w48221, w48222, w48223, w48224, w48225, w48226, w48227, w48228, w48229, w48230, w48231, w48232, w48233, w48234, w48235, w48236, w48237, w48238, w48239, w48240, w48241, w48242, w48243, w48244, w48245, w48246, w48247, w48248, w48249, w48250, w48251, w48252, w48253, w48254, w48255, w48256, w48257, w48258, w48259, w48260, w48261, w48262, w48263, w48264, w48265, w48266, w48267, w48268, w48269, w48270, w48271, w48272, w48273, w48274, w48275, w48276, w48277, w48278, w48279, w48280, w48281, w48282, w48283, w48284, w48285, w48286, w48287, w48288, w48289, w48290, w48291, w48292, w48293, w48294, w48295, w48296, w48297, w48298, w48299, w48300, w48301, w48302, w48303, w48304, w48305, w48306, w48307, w48308, w48309, w48310, w48311, w48312, w48313, w48314, w48315, w48316, w48317, w48318, w48319, w48320, w48321, w48322, w48323, w48324, w48325, w48326, w48327, w48328, w48329, w48330, w48331, w48332, w48333, w48334, w48335, w48336, w48337, w48338, w48339, w48340, w48341, w48342, w48343, w48344, w48345, w48346, w48347, w48348, w48349, w48350, w48351, w48352, w48353, w48354, w48355, w48356, w48357, w48358, w48359, w48360, w48361, w48362, w48363, w48364, w48365, w48366, w48367, w48368, w48369, w48370, w48371, w48372, w48373, w48374, w48375, w48376, w48377, w48378, w48379, w48380, w48381, w48382, w48383, w48384, w48385, w48386, w48387, w48388, w48389, w48390, w48391, w48392, w48393, w48394, w48395, w48396, w48397, w48398, w48399, w48400, w48401, w48402, w48403, w48404, w48405, w48406, w48407, w48408, w48409, w48410, w48411, w48412, w48413, w48414, w48415, w48416, w48417, w48418, w48419, w48420, w48421, w48422, w48423, w48424, w48425, w48426, w48427, w48428, w48429, w48430, w48431, w48432, w48433, w48434, w48435, w48436, w48437, w48438, w48439, w48440, w48441, w48442, w48443, w48444, w48445, w48446, w48447, w48448, w48449, w48450, w48451, w48452, w48453, w48454, w48455, w48456, w48457, w48458, w48459, w48460, w48461, w48462, w48463, w48464, w48465, w48466, w48467, w48468, w48469, w48470, w48471, w48472, w48473, w48474, w48475, w48476, w48477, w48478, w48479, w48480, w48481, w48482, w48483, w48484, w48485, w48486, w48487, w48488, w48489, w48490, w48491, w48492, w48493, w48494, w48495, w48496, w48497, w48498, w48499, w48500, w48501, w48502, w48503, w48504, w48505, w48506, w48507, w48508, w48509, w48510, w48511, w48512, w48513, w48514, w48515, w48516, w48517, w48518, w48519, w48520, w48521, w48522, w48523, w48524, w48525, w48526, w48527, w48528, w48529, w48530, w48531, w48532, w48533, w48534, w48535, w48536, w48537, w48538, w48539, w48540, w48541, w48542, w48543, w48544, w48545, w48546, w48547, w48548, w48549, w48550, w48551, w48552, w48553, w48554, w48555, w48556, w48557, w48558, w48559, w48560, w48561, w48562, w48563, w48564, w48565, w48566, w48567, w48568, w48569, w48570, w48571, w48572, w48573, w48574, w48575, w48576, w48577, w48578, w48579, w48580, w48581, w48582, w48583, w48584, w48585, w48586, w48587, w48588, w48589, w48590, w48591, w48592, w48593, w48594, w48595, w48596, w48597, w48598, w48599, w48600, w48601, w48602, w48603, w48604, w48605, w48606, w48607, w48608, w48609, w48610, w48611, w48612, w48613, w48614, w48615, w48616, w48617, w48618, w48619, w48620, w48621, w48622, w48623, w48624, w48625, w48626, w48627, w48628, w48629, w48630, w48631, w48632, w48633, w48634, w48635, w48636, w48637, w48638, w48639, w48640, w48641, w48642, w48643, w48644, w48645, w48646, w48647, w48648, w48649, w48650, w48651, w48652, w48653, w48654, w48655, w48656, w48657, w48658, w48659, w48660, w48661, w48662, w48663, w48664, w48665, w48666, w48667, w48668, w48669, w48670, w48671, w48672, w48673, w48674, w48675, w48676, w48677, w48678, w48679, w48680, w48681, w48682, w48683, w48684, w48685, w48686, w48687, w48688, w48689, w48690, w48691, w48692, w48693, w48694, w48695, w48696, w48697, w48698, w48699, w48700, w48701, w48702, w48703, w48704, w48705, w48706, w48707, w48708, w48709, w48710, w48711, w48712, w48713, w48714, w48715, w48716, w48717, w48718, w48719, w48720, w48721, w48722, w48723, w48724, w48725, w48726, w48727, w48728, w48729, w48730, w48731, w48732, w48733, w48734, w48735, w48736, w48737, w48738, w48739, w48740, w48741, w48742, w48743, w48744, w48745, w48746, w48747, w48748, w48749, w48750, w48751, w48752, w48753, w48754, w48755, w48756, w48757, w48758, w48759, w48760, w48761, w48762, w48763, w48764, w48765, w48766, w48767, w48768, w48769, w48770, w48771, w48772, w48773, w48774, w48775, w48776, w48777, w48778, w48779, w48780, w48781, w48782, w48783, w48784, w48785, w48786, w48787, w48788, w48789, w48790, w48791, w48792, w48793, w48794, w48795, w48796, w48797, w48798, w48799, w48800, w48801, w48802, w48803, w48804, w48805, w48806, w48807, w48808, w48809, w48810, w48811, w48812, w48813, w48814, w48815, w48816, w48817, w48818, w48819, w48820, w48821, w48822, w48823, w48824, w48825, w48826, w48827, w48828, w48829, w48830, w48831, w48832, w48833, w48834, w48835, w48836, w48837, w48838, w48839, w48840, w48841, w48842, w48843, w48844, w48845, w48846, w48847, w48848, w48849, w48850, w48851, w48852, w48853, w48854, w48855, w48856, w48857, w48858, w48859, w48860, w48861, w48862, w48863, w48864, w48865, w48866, w48867, w48868, w48869, w48870, w48871, w48872, w48873, w48874, w48875, w48876, w48877, w48878, w48879, w48880, w48881, w48882, w48883, w48884, w48885, w48886, w48887, w48888, w48889, w48890, w48891, w48892, w48893, w48894, w48895, w48896, w48897, w48898, w48899, w48900, w48901, w48902, w48903, w48904, w48905, w48906, w48907, w48908, w48909, w48910, w48911, w48912, w48913, w48914, w48915, w48916, w48917, w48918, w48919, w48920, w48921, w48922, w48923, w48924, w48925, w48926, w48927, w48928, w48929, w48930, w48931, w48932, w48933, w48934, w48935, w48936, w48937, w48938, w48939, w48940, w48941, w48942, w48943, w48944, w48945, w48946, w48947, w48948, w48949, w48950, w48951, w48952, w48953, w48954, w48955, w48956, w48957, w48958, w48959, w48960, w48961, w48962, w48963, w48964, w48965, w48966, w48967, w48968, w48969, w48970, w48971, w48972, w48973, w48974, w48975, w48976, w48977, w48978, w48979, w48980, w48981, w48982, w48983, w48984, w48985, w48986, w48987, w48988, w48989, w48990, w48991, w48992, w48993, w48994, w48995, w48996, w48997, w48998, w48999, w49000, w49001, w49002, w49003, w49004, w49005, w49006, w49007, w49008, w49009, w49010, w49011, w49012, w49013, w49014, w49015, w49016, w49017, w49018, w49019, w49020, w49021, w49022, w49023, w49024, w49025, w49026, w49027, w49028, w49029, w49030, w49031, w49032, w49033, w49034, w49035, w49036, w49037, w49038, w49039, w49040, w49041, w49042, w49043, w49044, w49045, w49046, w49047, w49048, w49049, w49050, w49051, w49052, w49053, w49054, w49055, w49056, w49057, w49058, w49059, w49060, w49061, w49062, w49063, w49064, w49065, w49066, w49067, w49068, w49069, w49070, w49071, w49072, w49073, w49074, w49075, w49076, w49077, w49078, w49079, w49080, w49081, w49082, w49083, w49084, w49085, w49086, w49087, w49088, w49089, w49090, w49091, w49092, w49093, w49094, w49095, w49096, w49097, w49098, w49099, w49100, w49101, w49102, w49103, w49104, w49105, w49106, w49107, w49108, w49109, w49110, w49111, w49112, w49113, w49114, w49115, w49116, w49117, w49118, w49119, w49120, w49121, w49122, w49123, w49124, w49125, w49126, w49127, w49128, w49129, w49130, w49131, w49132, w49133, w49134, w49135, w49136, w49137, w49138, w49139, w49140, w49141, w49142, w49143, w49144, w49145, w49146, w49147, w49148, w49149, w49150, w49151, w49152, w49153, w49154, w49155, w49156, w49157, w49158, w49159, w49160, w49161, w49162, w49163, w49164, w49165, w49166, w49167, w49168, w49169, w49170, w49171, w49172, w49173, w49174, w49175, w49176, w49177, w49178, w49179, w49180, w49181, w49182, w49183, w49184, w49185, w49186, w49187, w49188, w49189, w49190, w49191, w49192, w49193, w49194, w49195, w49196, w49197, w49198, w49199, w49200, w49201, w49202, w49203, w49204, w49205, w49206, w49207, w49208, w49209, w49210, w49211, w49212, w49213, w49214, w49215, w49216, w49217, w49218, w49219, w49220, w49221, w49222, w49223, w49224, w49225, w49226, w49227, w49228, w49229, w49230, w49231, w49232, w49233, w49234, w49235, w49236, w49237, w49238, w49239, w49240, w49241, w49242, w49243, w49244, w49245, w49246, w49247, w49248, w49249, w49250, w49251, w49252, w49253, w49254, w49255, w49256, w49257, w49258, w49259, w49260, w49261, w49262, w49263, w49264, w49265, w49266, w49267, w49268, w49269, w49270, w49271, w49272, w49273, w49274, w49275, w49276, w49277, w49278, w49279, w49280, w49281, w49282, w49283, w49284, w49285, w49286, w49287, w49288, w49289, w49290, w49291, w49292, w49293, w49294, w49295, w49296, w49297, w49298, w49299, w49300, w49301, w49302, w49303, w49304, w49305, w49306, w49307, w49308, w49309, w49310, w49311, w49312, w49313, w49314, w49315, w49316, w49317, w49318, w49319, w49320, w49321, w49322, w49323, w49324, w49325, w49326, w49327, w49328, w49329, w49330, w49331, w49332, w49333, w49334, w49335, w49336, w49337, w49338, w49339, w49340, w49341, w49342, w49343, w49344, w49345, w49346, w49347, w49348, w49349, w49350, w49351, w49352, w49353, w49354, w49355, w49356, w49357, w49358, w49359, w49360, w49361, w49362, w49363, w49364, w49365, w49366, w49367, w49368, w49369, w49370, w49371, w49372, w49373, w49374, w49375, w49376, w49377, w49378, w49379, w49380, w49381, w49382, w49383, w49384, w49385, w49386, w49387, w49388, w49389, w49390, w49391, w49392, w49393, w49394, w49395, w49396, w49397, w49398, w49399, w49400, w49401, w49402, w49403, w49404, w49405, w49406, w49407, w49408, w49409, w49410, w49411, w49412, w49413, w49414, w49415, w49416, w49417, w49418, w49419, w49420, w49421, w49422, w49423, w49424, w49425, w49426, w49427, w49428, w49429, w49430, w49431, w49432, w49433, w49434, w49435, w49436, w49437, w49438, w49439, w49440, w49441, w49442, w49443, w49444, w49445, w49446, w49447, w49448, w49449, w49450, w49451, w49452, w49453, w49454, w49455, w49456, w49457, w49458, w49459, w49460, w49461, w49462, w49463, w49464, w49465, w49466, w49467, w49468, w49469, w49470, w49471, w49472, w49473, w49474, w49475, w49476, w49477, w49478, w49479, w49480, w49481, w49482, w49483, w49484, w49485, w49486, w49487, w49488, w49489, w49490, w49491, w49492, w49493, w49494, w49495, w49496, w49497, w49498, w49499, w49500, w49501, w49502, w49503, w49504, w49505, w49506, w49507, w49508, w49509, w49510, w49511, w49512, w49513, w49514, w49515, w49516, w49517, w49518, w49519, w49520, w49521, w49522, w49523, w49524, w49525, w49526, w49527, w49528, w49529, w49530, w49531, w49532, w49533, w49534, w49535, w49536, w49537, w49538, w49539, w49540, w49541, w49542, w49543, w49544, w49545, w49546, w49547, w49548, w49549, w49550, w49551, w49552, w49553, w49554, w49555, w49556, w49557, w49558, w49559, w49560, w49561, w49562, w49563, w49564, w49565, w49566, w49567, w49568, w49569, w49570, w49571, w49572, w49573, w49574, w49575, w49576, w49577, w49578, w49579, w49580, w49581, w49582, w49583, w49584, w49585, w49586, w49587, w49588, w49589, w49590, w49591, w49592, w49593, w49594, w49595, w49596, w49597, w49598, w49599, w49600, w49601, w49602, w49603, w49604, w49605, w49606, w49607, w49608, w49609, w49610, w49611, w49612, w49613, w49614, w49615, w49616, w49617, w49618, w49619, w49620, w49621, w49622, w49623, w49624, w49625, w49626, w49627, w49628, w49629, w49630, w49631, w49632, w49633, w49634, w49635, w49636, w49637, w49638, w49639, w49640, w49641, w49642, w49643, w49644, w49645, w49646, w49647, w49648, w49649, w49650, w49651, w49652, w49653, w49654, w49655, w49656, w49657, w49658, w49659, w49660, w49661, w49662, w49663, w49664, w49665, w49666, w49667, w49668, w49669, w49670, w49671, w49672, w49673, w49674, w49675, w49676, w49677, w49678, w49679, w49680, w49681, w49682, w49683, w49684, w49685, w49686, w49687, w49688, w49689, w49690, w49691, w49692, w49693, w49694, w49695, w49696, w49697, w49698, w49699, w49700, w49701, w49702, w49703, w49704, w49705, w49706, w49707, w49708, w49709, w49710, w49711, w49712, w49713, w49714, w49715, w49716, w49717, w49718, w49719, w49720, w49721, w49722, w49723, w49724, w49725, w49726, w49727, w49728, w49729, w49730, w49731, w49732, w49733, w49734, w49735, w49736, w49737, w49738, w49739, w49740, w49741, w49742, w49743, w49744, w49745, w49746, w49747, w49748, w49749, w49750, w49751, w49752, w49753, w49754, w49755, w49756, w49757, w49758, w49759, w49760, w49761, w49762, w49763, w49764, w49765, w49766, w49767, w49768, w49769, w49770, w49771, w49772, w49773, w49774, w49775, w49776, w49777, w49778, w49779, w49780, w49781, w49782, w49783, w49784, w49785, w49786, w49787, w49788, w49789, w49790, w49791, w49792, w49793, w49794, w49795, w49796, w49797, w49798, w49799, w49800, w49801, w49802, w49803, w49804, w49805, w49806, w49807, w49808, w49809, w49810, w49811, w49812, w49813, w49814, w49815, w49816, w49817, w49818, w49819, w49820, w49821, w49822, w49823, w49824, w49825, w49826, w49827, w49828, w49829, w49830, w49831, w49832, w49833, w49834, w49835, w49836, w49837, w49838, w49839, w49840, w49841, w49842, w49843, w49844, w49845, w49846, w49847, w49848, w49849, w49850, w49851, w49852, w49853, w49854, w49855, w49856, w49857, w49858, w49859, w49860, w49861, w49862, w49863, w49864, w49865, w49866, w49867, w49868, w49869, w49870, w49871, w49872, w49873, w49874, w49875, w49876, w49877, w49878, w49879, w49880, w49881, w49882, w49883, w49884, w49885, w49886, w49887, w49888, w49889, w49890, w49891, w49892, w49893, w49894, w49895, w49896, w49897, w49898, w49899, w49900, w49901, w49902, w49903, w49904, w49905, w49906, w49907, w49908, w49909, w49910, w49911, w49912, w49913, w49914, w49915, w49916, w49917, w49918, w49919, w49920, w49921, w49922, w49923, w49924, w49925, w49926, w49927, w49928, w49929, w49930, w49931, w49932, w49933, w49934, w49935, w49936, w49937, w49938, w49939, w49940, w49941, w49942, w49943, w49944, w49945, w49946, w49947, w49948, w49949, w49950, w49951, w49952, w49953, w49954, w49955, w49956, w49957, w49958, w49959, w49960, w49961, w49962, w49963, w49964, w49965, w49966, w49967, w49968, w49969, w49970, w49971, w49972, w49973, w49974, w49975, w49976, w49977, w49978, w49979, w49980, w49981, w49982, w49983, w49984, w49985, w49986, w49987, w49988, w49989, w49990, w49991, w49992, w49993, w49994, w49995, w49996, w49997, w49998, w49999, w50000, w50001, w50002, w50003, w50004, w50005, w50006, w50007, w50008, w50009, w50010, w50011, w50012, w50013, w50014, w50015, w50016, w50017, w50018, w50019, w50020, w50021, w50022, w50023, w50024, w50025, w50026, w50027, w50028, w50029, w50030, w50031, w50032, w50033, w50034, w50035, w50036, w50037, w50038, w50039, w50040, w50041, w50042, w50043, w50044, w50045, w50046, w50047, w50048, w50049, w50050, w50051, w50052, w50053, w50054, w50055, w50056, w50057, w50058, w50059, w50060, w50061, w50062, w50063, w50064, w50065, w50066, w50067, w50068, w50069, w50070, w50071, w50072, w50073, w50074, w50075, w50076, w50077, w50078, w50079, w50080, w50081, w50082, w50083, w50084, w50085, w50086, w50087, w50088, w50089, w50090, w50091, w50092, w50093, w50094, w50095, w50096, w50097, w50098, w50099, w50100, w50101, w50102, w50103, w50104, w50105, w50106, w50107, w50108, w50109, w50110, w50111, w50112, w50113, w50114, w50115, w50116, w50117, w50118, w50119, w50120, w50121, w50122, w50123, w50124, w50125, w50126, w50127, w50128, w50129, w50130, w50131, w50132, w50133, w50134, w50135, w50136, w50137, w50138, w50139, w50140, w50141, w50142, w50143, w50144, w50145, w50146, w50147, w50148, w50149, w50150, w50151, w50152, w50153, w50154, w50155, w50156, w50157, w50158, w50159, w50160, w50161, w50162, w50163, w50164, w50165, w50166, w50167, w50168, w50169, w50170, w50171, w50172, w50173, w50174, w50175, w50176, w50177, w50178, w50179, w50180, w50181, w50182, w50183, w50184, w50185, w50186, w50187, w50188, w50189, w50190, w50191, w50192, w50193, w50194, w50195, w50196, w50197, w50198, w50199, w50200, w50201, w50202, w50203, w50204, w50205, w50206, w50207, w50208, w50209, w50210, w50211, w50212, w50213, w50214, w50215, w50216, w50217, w50218, w50219, w50220, w50221, w50222, w50223, w50224, w50225, w50226, w50227, w50228, w50229, w50230, w50231, w50232, w50233, w50234, w50235, w50236, w50237, w50238, w50239, w50240, w50241, w50242, w50243, w50244, w50245, w50246, w50247, w50248, w50249, w50250, w50251, w50252, w50253, w50254, w50255, w50256, w50257, w50258, w50259, w50260, w50261, w50262, w50263, w50264, w50265, w50266, w50267, w50268, w50269, w50270, w50271, w50272, w50273, w50274, w50275, w50276, w50277, w50278, w50279, w50280, w50281, w50282, w50283, w50284, w50285, w50286, w50287, w50288, w50289, w50290, w50291, w50292, w50293, w50294, w50295, w50296, w50297, w50298, w50299, w50300, w50301, w50302, w50303, w50304, w50305, w50306, w50307, w50308, w50309, w50310, w50311, w50312, w50313, w50314, w50315, w50316, w50317, w50318, w50319, w50320, w50321, w50322, w50323, w50324, w50325, w50326, w50327, w50328, w50329, w50330, w50331, w50332, w50333, w50334, w50335, w50336, w50337, w50338, w50339, w50340, w50341, w50342, w50343, w50344, w50345, w50346, w50347, w50348, w50349, w50350, w50351, w50352, w50353, w50354, w50355, w50356, w50357, w50358, w50359, w50360, w50361, w50362, w50363, w50364, w50365, w50366, w50367, w50368, w50369, w50370, w50371, w50372, w50373, w50374, w50375, w50376, w50377, w50378, w50379, w50380, w50381, w50382, w50383, w50384, w50385, w50386, w50387, w50388, w50389, w50390, w50391, w50392, w50393, w50394, w50395, w50396, w50397, w50398, w50399, w50400, w50401, w50402, w50403, w50404, w50405, w50406, w50407, w50408, w50409, w50410, w50411, w50412, w50413, w50414, w50415, w50416, w50417, w50418, w50419, w50420, w50421, w50422, w50423, w50424, w50425, w50426, w50427, w50428, w50429, w50430, w50431, w50432, w50433, w50434, w50435, w50436, w50437, w50438, w50439, w50440, w50441, w50442, w50443, w50444, w50445, w50446, w50447, w50448, w50449, w50450, w50451, w50452, w50453, w50454, w50455, w50456, w50457, w50458, w50459, w50460, w50461, w50462, w50463, w50464, w50465, w50466, w50467, w50468, w50469, w50470, w50471, w50472, w50473, w50474, w50475, w50476, w50477, w50478, w50479, w50480, w50481, w50482, w50483, w50484, w50485, w50486, w50487, w50488, w50489, w50490, w50491, w50492, w50493, w50494, w50495, w50496, w50497, w50498, w50499, w50500, w50501, w50502, w50503, w50504, w50505, w50506, w50507, w50508, w50509, w50510, w50511, w50512, w50513, w50514, w50515, w50516, w50517, w50518, w50519, w50520, w50521, w50522, w50523, w50524, w50525, w50526, w50527, w50528, w50529, w50530, w50531, w50532, w50533, w50534, w50535, w50536, w50537, w50538, w50539, w50540, w50541, w50542, w50543, w50544, w50545, w50546, w50547, w50548, w50549, w50550, w50551, w50552, w50553, w50554, w50555, w50556, w50557, w50558, w50559, w50560, w50561, w50562, w50563, w50564, w50565, w50566, w50567, w50568, w50569, w50570, w50571, w50572, w50573, w50574, w50575, w50576, w50577, w50578, w50579, w50580, w50581, w50582, w50583, w50584, w50585, w50586, w50587, w50588, w50589, w50590, w50591, w50592, w50593, w50594, w50595, w50596, w50597, w50598, w50599, w50600, w50601, w50602, w50603, w50604, w50605, w50606, w50607, w50608, w50609, w50610, w50611, w50612, w50613, w50614, w50615, w50616, w50617, w50618, w50619, w50620, w50621, w50622, w50623, w50624, w50625, w50626, w50627, w50628, w50629, w50630, w50631, w50632, w50633, w50634, w50635, w50636, w50637, w50638, w50639, w50640, w50641, w50642, w50643, w50644, w50645, w50646, w50647, w50648, w50649, w50650, w50651, w50652, w50653, w50654, w50655, w50656, w50657, w50658, w50659, w50660, w50661, w50662, w50663, w50664, w50665, w50666, w50667, w50668, w50669, w50670, w50671, w50672, w50673, w50674, w50675, w50676, w50677, w50678, w50679, w50680, w50681, w50682, w50683, w50684, w50685, w50686, w50687, w50688, w50689, w50690, w50691, w50692, w50693, w50694, w50695, w50696, w50697, w50698, w50699, w50700, w50701, w50702, w50703, w50704, w50705, w50706, w50707, w50708, w50709, w50710, w50711, w50712, w50713, w50714, w50715, w50716, w50717, w50718, w50719, w50720, w50721, w50722, w50723, w50724, w50725, w50726, w50727, w50728, w50729, w50730, w50731, w50732, w50733, w50734, w50735, w50736, w50737, w50738, w50739, w50740, w50741, w50742, w50743, w50744, w50745, w50746, w50747, w50748, w50749, w50750, w50751, w50752, w50753, w50754, w50755, w50756, w50757, w50758, w50759, w50760, w50761, w50762, w50763, w50764, w50765, w50766, w50767, w50768, w50769, w50770, w50771, w50772, w50773, w50774, w50775, w50776, w50777, w50778, w50779, w50780, w50781, w50782, w50783, w50784, w50785, w50786, w50787, w50788, w50789, w50790, w50791, w50792, w50793, w50794, w50795, w50796, w50797, w50798, w50799, w50800, w50801, w50802, w50803, w50804, w50805, w50806, w50807, w50808, w50809, w50810, w50811, w50812, w50813, w50814, w50815, w50816, w50817, w50818, w50819, w50820, w50821, w50822, w50823, w50824, w50825, w50826, w50827, w50828, w50829, w50830, w50831, w50832, w50833, w50834, w50835, w50836, w50837, w50838, w50839, w50840, w50841, w50842, w50843, w50844, w50845, w50846, w50847, w50848, w50849, w50850, w50851, w50852, w50853, w50854, w50855, w50856, w50857, w50858, w50859, w50860, w50861, w50862, w50863, w50864, w50865, w50866, w50867, w50868, w50869, w50870, w50871, w50872, w50873, w50874, w50875, w50876, w50877, w50878, w50879, w50880, w50881, w50882, w50883, w50884, w50885, w50886, w50887, w50888, w50889, w50890, w50891, w50892, w50893, w50894, w50895, w50896, w50897, w50898, w50899, w50900, w50901, w50902, w50903, w50904, w50905, w50906, w50907, w50908, w50909, w50910, w50911, w50912, w50913, w50914, w50915, w50916, w50917, w50918, w50919, w50920, w50921;

	assign w47765 = w383 ^ w255;
	assign w47766 = w382 ^ w254;
	assign w47767 = w381 ^ w253;
	assign w47768 = w380 ^ w252;
	assign w47769 = w379 ^ w251;
	assign w47770 = w378 ^ w250;
	assign w47771 = w377 ^ w249;
	assign w47772 = w376 ^ w248;
	assign w47773 = w375 ^ w247;
	assign w47774 = w374 ^ w246;
	assign w47775 = w373 ^ w245;
	assign w47776 = w372 ^ w244;
	assign w47777 = w371 ^ w243;
	assign w47778 = w370 ^ w242;
	assign w47779 = w369 ^ w241;
	assign w47780 = w368 ^ w240;
	assign w47781 = w367 ^ w239;
	assign w47782 = w366 ^ w238;
	assign w47783 = w365 ^ w237;
	assign w47784 = w364 ^ w236;
	assign w47785 = w363 ^ w235;
	assign w47786 = w362 ^ w234;
	assign w47787 = w361 ^ w233;
	assign w47788 = w360 ^ w232;
	assign w47789 = w359 ^ w231;
	assign w47790 = w358 ^ w230;
	assign w47791 = w357 ^ w229;
	assign w47792 = w356 ^ w228;
	assign w47793 = w355 ^ w227;
	assign w47794 = w354 ^ w226;
	assign w47795 = w353 ^ w225;
	assign w47796 = w352 ^ w224;
	assign w47797 = w351 ^ w223;
	assign w47798 = w350 ^ w222;
	assign w47799 = w349 ^ w221;
	assign w47800 = w348 ^ w220;
	assign w47801 = w347 ^ w219;
	assign w47802 = w346 ^ w218;
	assign w47803 = w345 ^ w217;
	assign w47804 = w344 ^ w216;
	assign w47805 = w343 ^ w215;
	assign w47806 = w342 ^ w214;
	assign w47807 = w341 ^ w213;
	assign w47808 = w340 ^ w212;
	assign w47809 = w339 ^ w211;
	assign w47810 = w338 ^ w210;
	assign w47811 = w337 ^ w209;
	assign w47812 = w336 ^ w208;
	assign w47813 = w335 ^ w207;
	assign w47814 = w334 ^ w206;
	assign w47815 = w333 ^ w205;
	assign w47816 = w332 ^ w204;
	assign w47817 = w331 ^ w203;
	assign w47818 = w330 ^ w202;
	assign w47819 = w329 ^ w201;
	assign w47820 = w328 ^ w200;
	assign w47821 = w327 ^ w199;
	assign w47822 = w326 ^ w198;
	assign w47823 = w325 ^ w197;
	assign w47824 = w324 ^ w196;
	assign w47825 = w323 ^ w195;
	assign w47826 = w322 ^ w194;
	assign w47827 = w321 ^ w193;
	assign w47828 = w320 ^ w192;
	assign w47829 = w319 ^ w191;
	assign w47830 = w318 ^ w190;
	assign w47831 = w317 ^ w189;
	assign w47832 = w316 ^ w188;
	assign w47833 = w315 ^ w187;
	assign w47834 = w314 ^ w186;
	assign w47835 = w313 ^ w185;
	assign w47836 = w312 ^ w184;
	assign w47837 = w311 ^ w183;
	assign w47838 = w310 ^ w182;
	assign w47839 = w309 ^ w181;
	assign w47840 = w308 ^ w180;
	assign w47841 = w307 ^ w179;
	assign w47842 = w306 ^ w178;
	assign w47843 = w305 ^ w177;
	assign w47844 = w304 ^ w176;
	assign w47845 = w303 ^ w175;
	assign w47846 = w302 ^ w174;
	assign w47847 = w301 ^ w173;
	assign w47848 = w300 ^ w172;
	assign w47849 = w299 ^ w171;
	assign w47850 = w298 ^ w170;
	assign w47851 = w297 ^ w169;
	assign w47852 = w296 ^ w168;
	assign w47853 = w295 ^ w167;
	assign w47854 = w294 ^ w166;
	assign w47855 = w293 ^ w165;
	assign w47856 = w292 ^ w164;
	assign w47857 = w291 ^ w163;
	assign w47858 = w290 ^ w162;
	assign w47859 = w289 ^ w161;
	assign w47860 = w288 ^ w160;
	assign w47861 = w287 ^ w159;
	assign w47862 = w286 ^ w158;
	assign w47863 = w285 ^ w157;
	assign w47864 = w284 ^ w156;
	assign w47865 = w283 ^ w155;
	assign w47866 = w282 ^ w154;
	assign w47867 = w281 ^ w153;
	assign w47868 = w280 ^ w152;
	assign w47869 = w279 ^ w151;
	assign w47870 = w278 ^ w150;
	assign w47871 = w277 ^ w149;
	assign w47872 = w276 ^ w148;
	assign w47873 = w275 ^ w147;
	assign w47874 = w274 ^ w146;
	assign w47875 = w273 ^ w145;
	assign w47876 = w272 ^ w144;
	assign w47877 = w271 ^ w143;
	assign w47878 = w270 ^ w142;
	assign w47879 = w269 ^ w141;
	assign w47880 = w268 ^ w140;
	assign w47881 = w267 ^ w139;
	assign w47882 = w266 ^ w138;
	assign w47883 = w265 ^ w137;
	assign w47884 = w264 ^ w136;
	assign w47885 = w263 ^ w135;
	assign w47886 = w262 ^ w134;
	assign w47887 = w261 ^ w133;
	assign w47888 = w260 ^ w132;
	assign w47889 = w259 ^ w131;
	assign w47890 = w258 ^ w130;
	assign w47891 = w257 ^ w129;
	assign w47892 = w256 ^ w128;
	assign w3547 = w17 ^ w19;
	assign w3546 = w21 ^ w23;
	assign w3545 = w18 ^ w3547;
	assign w3639 = w22 ^ w3545;
	assign w3636 = w21 ^ w3545;
	assign w3544 = w20 ^ w22;
	assign w3540 = w16 ^ w22;
	assign w3638 = w3540 ^ w3545;
	assign w3650 = w20 ^ w23;
	assign w3645 = w3546 ^ w3540;
	assign w3642 = w3547 ^ w3650;
	assign w3641 = w16 ^ w3642;
	assign w3529 = w17 ^ w18;
	assign w3643 = w3529 ^ w3645;
	assign w3646 = w3650 ^ w3529;
	assign w3652 = w18 ^ w20;
	assign w3637 = w3546 ^ w3652;
	assign w3648 = w21 ^ w3540;
	assign w3644 = w17 ^ w3648;
	assign w3570 = w19 ^ w18;
	assign w3584 = w3544 ^ w3546;
	assign w3640 = w3547 ^ w3584;
	assign w3585 = w3544 ^ w21;
	assign w3647 = w16 ^ w3585;
	assign w3651 = w23 ^ w17;
	assign w3649 = w23 ^ w18;
	assign w3635 = w3642 & w3646;
	assign w3541 = w3635 ^ w3544;
	assign w3634 = w3643 & w3641;
	assign w3633 = w3647 & w16;
	assign w3632 = w3651 & w3636;
	assign w3542 = w3632 ^ w3546;
	assign w3631 = w3648 & w3644;
	assign w3630 = w3645 & w3638;
	assign w3629 = w3650 & w3639;
	assign w3543 = w3629 ^ w3545;
	assign w3537 = w3541 ^ w3543;
	assign w3531 = w23 ^ w3537;
	assign w3628 = w3652 & w3637;
	assign w3536 = w3628 ^ w3634;
	assign w3626 = w3536 ^ w3531;
	assign w3571 = w3628 ^ w3629;
	assign w3523 = w3571 ^ w3570;
	assign w3524 = w3523 ^ w3542;
	assign w3625 = w3631 ^ w3524;
	assign w3627 = w3649 & w3640;
	assign w3622 = w3626 & w3625;
	assign w3695 = w9 ^ w11;
	assign w3696 = w13 ^ w15;
	assign w3697 = w10 ^ w3695;
	assign w3773 = w14 ^ w3697;
	assign w3770 = w13 ^ w3697;
	assign w3698 = w12 ^ w14;
	assign w3702 = w8 ^ w14;
	assign w3772 = w3702 ^ w3697;
	assign w3784 = w12 ^ w15;
	assign w3779 = w3696 ^ w3702;
	assign w3776 = w3695 ^ w3784;
	assign w3775 = w8 ^ w3776;
	assign w3712 = w9 ^ w10;
	assign w3777 = w3712 ^ w3779;
	assign w3780 = w3784 ^ w3712;
	assign w3786 = w10 ^ w12;
	assign w3771 = w3696 ^ w3786;
	assign w3782 = w13 ^ w3702;
	assign w3778 = w9 ^ w3782;
	assign w3672 = w11 ^ w10;
	assign w3658 = w3698 ^ w3696;
	assign w3774 = w3695 ^ w3658;
	assign w3657 = w3698 ^ w13;
	assign w3781 = w8 ^ w3657;
	assign w3785 = w15 ^ w9;
	assign w3783 = w15 ^ w10;
	assign w3769 = w3776 & w3780;
	assign w3701 = w3769 ^ w3698;
	assign w3768 = w3777 & w3775;
	assign w3767 = w3781 & w8;
	assign w3766 = w3785 & w3770;
	assign w3700 = w3766 ^ w3696;
	assign w3765 = w3782 & w3778;
	assign w3764 = w3779 & w3772;
	assign w3763 = w3784 & w3773;
	assign w3699 = w3763 ^ w3697;
	assign w3705 = w3701 ^ w3699;
	assign w3710 = w15 ^ w3705;
	assign w3762 = w3786 & w3771;
	assign w3719 = w3762 ^ w3768;
	assign w3760 = w3719 ^ w3710;
	assign w3671 = w3762 ^ w3763;
	assign w3718 = w3671 ^ w3672;
	assign w3717 = w3718 ^ w3700;
	assign w3759 = w3765 ^ w3717;
	assign w3761 = w3783 & w3774;
	assign w3756 = w3760 & w3759;
	assign w3829 = w1 ^ w3;
	assign w3830 = w5 ^ w7;
	assign w3831 = w2 ^ w3829;
	assign w3907 = w6 ^ w3831;
	assign w3904 = w5 ^ w3831;
	assign w3832 = w4 ^ w6;
	assign w3836 = w0 ^ w6;
	assign w3906 = w3836 ^ w3831;
	assign w3918 = w4 ^ w7;
	assign w3913 = w3830 ^ w3836;
	assign w3910 = w3829 ^ w3918;
	assign w3909 = w0 ^ w3910;
	assign w3846 = w1 ^ w2;
	assign w3911 = w3846 ^ w3913;
	assign w3914 = w3918 ^ w3846;
	assign w3920 = w2 ^ w4;
	assign w3905 = w3830 ^ w3920;
	assign w3916 = w5 ^ w3836;
	assign w3912 = w1 ^ w3916;
	assign w3806 = w3 ^ w2;
	assign w3792 = w3832 ^ w3830;
	assign w3908 = w3829 ^ w3792;
	assign w3791 = w3832 ^ w5;
	assign w3915 = w0 ^ w3791;
	assign w3919 = w7 ^ w1;
	assign w3917 = w7 ^ w2;
	assign w3903 = w3910 & w3914;
	assign w3835 = w3903 ^ w3832;
	assign w3902 = w3911 & w3909;
	assign w3901 = w3915 & w0;
	assign w3900 = w3919 & w3904;
	assign w3834 = w3900 ^ w3830;
	assign w3899 = w3916 & w3912;
	assign w3898 = w3913 & w3906;
	assign w3897 = w3918 & w3907;
	assign w3833 = w3897 ^ w3831;
	assign w3839 = w3835 ^ w3833;
	assign w3844 = w7 ^ w3839;
	assign w3896 = w3920 & w3905;
	assign w3853 = w3896 ^ w3902;
	assign w3894 = w3853 ^ w3844;
	assign w3805 = w3896 ^ w3897;
	assign w3852 = w3805 ^ w3806;
	assign w3851 = w3852 ^ w3834;
	assign w3893 = w3899 ^ w3851;
	assign w3895 = w3917 & w3908;
	assign w3890 = w3894 & w3893;
	assign w3963 = w25 ^ w27;
	assign w3964 = w29 ^ w31;
	assign w3965 = w26 ^ w3963;
	assign w4041 = w30 ^ w3965;
	assign w4038 = w29 ^ w3965;
	assign w3966 = w28 ^ w30;
	assign w3970 = w24 ^ w30;
	assign w4040 = w3970 ^ w3965;
	assign w4052 = w28 ^ w31;
	assign w4047 = w3964 ^ w3970;
	assign w4044 = w3963 ^ w4052;
	assign w4043 = w24 ^ w4044;
	assign w3980 = w25 ^ w26;
	assign w4045 = w3980 ^ w4047;
	assign w4048 = w4052 ^ w3980;
	assign w4054 = w26 ^ w28;
	assign w4039 = w3964 ^ w4054;
	assign w4050 = w29 ^ w3970;
	assign w4046 = w25 ^ w4050;
	assign w3940 = w27 ^ w26;
	assign w3926 = w3966 ^ w3964;
	assign w4042 = w3963 ^ w3926;
	assign w3925 = w3966 ^ w29;
	assign w4049 = w24 ^ w3925;
	assign w4053 = w31 ^ w25;
	assign w4051 = w31 ^ w26;
	assign w4037 = w4044 & w4048;
	assign w3969 = w4037 ^ w3966;
	assign w4036 = w4045 & w4043;
	assign w4035 = w4049 & w24;
	assign w4034 = w4053 & w4038;
	assign w3968 = w4034 ^ w3964;
	assign w4033 = w4050 & w4046;
	assign w4032 = w4047 & w4040;
	assign w4031 = w4052 & w4041;
	assign w3967 = w4031 ^ w3965;
	assign w3973 = w3969 ^ w3967;
	assign w3978 = w31 ^ w3973;
	assign w4030 = w4054 & w4039;
	assign w3987 = w4030 ^ w4036;
	assign w4028 = w3987 ^ w3978;
	assign w3939 = w4030 ^ w4031;
	assign w3986 = w3939 ^ w3940;
	assign w3985 = w3986 ^ w3968;
	assign w4027 = w4033 ^ w3985;
	assign w4029 = w4051 & w4042;
	assign w4024 = w4028 & w4027;
	assign w5172 = w47883 ^ w47881;
	assign w5173 = w47879 ^ w47877;
	assign w5174 = w47882 ^ w5172;
	assign w5250 = w47878 ^ w5174;
	assign w5247 = w47879 ^ w5174;
	assign w5175 = w47880 ^ w47878;
	assign w5179 = w47884 ^ w47878;
	assign w5249 = w5179 ^ w5174;
	assign w5261 = w47880 ^ w47877;
	assign w5256 = w5173 ^ w5179;
	assign w5253 = w5172 ^ w5261;
	assign w5252 = w47884 ^ w5253;
	assign w5189 = w47883 ^ w47882;
	assign w5254 = w5189 ^ w5256;
	assign w5257 = w5261 ^ w5189;
	assign w5263 = w47882 ^ w47880;
	assign w5248 = w5173 ^ w5263;
	assign w5259 = w47879 ^ w5179;
	assign w5255 = w47883 ^ w5259;
	assign w5149 = w47881 ^ w47882;
	assign w5135 = w5175 ^ w5173;
	assign w5251 = w5172 ^ w5135;
	assign w5134 = w5175 ^ w47879;
	assign w5258 = w47884 ^ w5134;
	assign w5262 = w47877 ^ w47883;
	assign w5260 = w47877 ^ w47882;
	assign w5246 = w5253 & w5257;
	assign w5178 = w5246 ^ w5175;
	assign w5245 = w5254 & w5252;
	assign w5244 = w5258 & w47884;
	assign w5243 = w5262 & w5247;
	assign w5177 = w5243 ^ w5173;
	assign w5242 = w5259 & w5255;
	assign w5241 = w5256 & w5249;
	assign w5240 = w5261 & w5250;
	assign w5176 = w5240 ^ w5174;
	assign w5182 = w5178 ^ w5176;
	assign w5187 = w47877 ^ w5182;
	assign w5239 = w5263 & w5248;
	assign w5196 = w5239 ^ w5245;
	assign w5237 = w5196 ^ w5187;
	assign w5148 = w5239 ^ w5240;
	assign w5195 = w5148 ^ w5149;
	assign w5194 = w5195 ^ w5177;
	assign w5236 = w5242 ^ w5194;
	assign w5238 = w5260 & w5251;
	assign w5233 = w5237 & w5236;
	assign w5306 = w47875 ^ w47873;
	assign w5307 = w47871 ^ w47869;
	assign w5308 = w47874 ^ w5306;
	assign w5384 = w47870 ^ w5308;
	assign w5381 = w47871 ^ w5308;
	assign w5309 = w47872 ^ w47870;
	assign w5313 = w47876 ^ w47870;
	assign w5383 = w5313 ^ w5308;
	assign w5395 = w47872 ^ w47869;
	assign w5390 = w5307 ^ w5313;
	assign w5387 = w5306 ^ w5395;
	assign w5386 = w47876 ^ w5387;
	assign w5323 = w47875 ^ w47874;
	assign w5388 = w5323 ^ w5390;
	assign w5391 = w5395 ^ w5323;
	assign w5397 = w47874 ^ w47872;
	assign w5382 = w5307 ^ w5397;
	assign w5393 = w47871 ^ w5313;
	assign w5389 = w47875 ^ w5393;
	assign w5283 = w47873 ^ w47874;
	assign w5269 = w5309 ^ w5307;
	assign w5385 = w5306 ^ w5269;
	assign w5268 = w5309 ^ w47871;
	assign w5392 = w47876 ^ w5268;
	assign w5396 = w47869 ^ w47875;
	assign w5394 = w47869 ^ w47874;
	assign w5380 = w5387 & w5391;
	assign w5312 = w5380 ^ w5309;
	assign w5379 = w5388 & w5386;
	assign w5378 = w5392 & w47876;
	assign w5377 = w5396 & w5381;
	assign w5311 = w5377 ^ w5307;
	assign w5376 = w5393 & w5389;
	assign w5375 = w5390 & w5383;
	assign w5374 = w5395 & w5384;
	assign w5310 = w5374 ^ w5308;
	assign w5316 = w5312 ^ w5310;
	assign w5321 = w47869 ^ w5316;
	assign w5373 = w5397 & w5382;
	assign w5330 = w5373 ^ w5379;
	assign w5371 = w5330 ^ w5321;
	assign w5282 = w5373 ^ w5374;
	assign w5329 = w5282 ^ w5283;
	assign w5328 = w5329 ^ w5311;
	assign w5370 = w5376 ^ w5328;
	assign w5372 = w5394 & w5385;
	assign w5367 = w5371 & w5370;
	assign w5440 = w47867 ^ w47865;
	assign w5441 = w47863 ^ w47861;
	assign w5442 = w47866 ^ w5440;
	assign w5518 = w47862 ^ w5442;
	assign w5515 = w47863 ^ w5442;
	assign w5443 = w47864 ^ w47862;
	assign w5447 = w47868 ^ w47862;
	assign w5517 = w5447 ^ w5442;
	assign w5529 = w47864 ^ w47861;
	assign w5524 = w5441 ^ w5447;
	assign w5521 = w5440 ^ w5529;
	assign w5520 = w47868 ^ w5521;
	assign w5457 = w47867 ^ w47866;
	assign w5522 = w5457 ^ w5524;
	assign w5525 = w5529 ^ w5457;
	assign w5531 = w47866 ^ w47864;
	assign w5516 = w5441 ^ w5531;
	assign w5527 = w47863 ^ w5447;
	assign w5523 = w47867 ^ w5527;
	assign w5417 = w47865 ^ w47866;
	assign w5403 = w5443 ^ w5441;
	assign w5519 = w5440 ^ w5403;
	assign w5402 = w5443 ^ w47863;
	assign w5526 = w47868 ^ w5402;
	assign w5530 = w47861 ^ w47867;
	assign w5528 = w47861 ^ w47866;
	assign w5514 = w5521 & w5525;
	assign w5446 = w5514 ^ w5443;
	assign w5513 = w5522 & w5520;
	assign w5512 = w5526 & w47868;
	assign w5511 = w5530 & w5515;
	assign w5445 = w5511 ^ w5441;
	assign w5510 = w5527 & w5523;
	assign w5509 = w5524 & w5517;
	assign w5508 = w5529 & w5518;
	assign w5444 = w5508 ^ w5442;
	assign w5450 = w5446 ^ w5444;
	assign w5455 = w47861 ^ w5450;
	assign w5507 = w5531 & w5516;
	assign w5464 = w5507 ^ w5513;
	assign w5505 = w5464 ^ w5455;
	assign w5416 = w5507 ^ w5508;
	assign w5463 = w5416 ^ w5417;
	assign w5462 = w5463 ^ w5445;
	assign w5504 = w5510 ^ w5462;
	assign w5506 = w5528 & w5519;
	assign w5501 = w5505 & w5504;
	assign w5574 = w47851 ^ w47849;
	assign w5575 = w47847 ^ w47845;
	assign w5576 = w47850 ^ w5574;
	assign w5652 = w47846 ^ w5576;
	assign w5649 = w47847 ^ w5576;
	assign w5577 = w47848 ^ w47846;
	assign w5581 = w47852 ^ w47846;
	assign w5651 = w5581 ^ w5576;
	assign w5663 = w47848 ^ w47845;
	assign w5658 = w5575 ^ w5581;
	assign w5655 = w5574 ^ w5663;
	assign w5654 = w47852 ^ w5655;
	assign w5591 = w47851 ^ w47850;
	assign w5656 = w5591 ^ w5658;
	assign w5659 = w5663 ^ w5591;
	assign w5665 = w47850 ^ w47848;
	assign w5650 = w5575 ^ w5665;
	assign w5661 = w47847 ^ w5581;
	assign w5657 = w47851 ^ w5661;
	assign w5551 = w47849 ^ w47850;
	assign w5537 = w5577 ^ w5575;
	assign w5653 = w5574 ^ w5537;
	assign w5536 = w5577 ^ w47847;
	assign w5660 = w47852 ^ w5536;
	assign w5664 = w47845 ^ w47851;
	assign w5662 = w47845 ^ w47850;
	assign w5648 = w5655 & w5659;
	assign w5580 = w5648 ^ w5577;
	assign w5647 = w5656 & w5654;
	assign w5646 = w5660 & w47852;
	assign w5645 = w5664 & w5649;
	assign w5579 = w5645 ^ w5575;
	assign w5644 = w5661 & w5657;
	assign w5643 = w5658 & w5651;
	assign w5642 = w5663 & w5652;
	assign w5578 = w5642 ^ w5576;
	assign w5584 = w5580 ^ w5578;
	assign w5589 = w47845 ^ w5584;
	assign w5641 = w5665 & w5650;
	assign w5598 = w5641 ^ w5647;
	assign w5639 = w5598 ^ w5589;
	assign w5550 = w5641 ^ w5642;
	assign w5597 = w5550 ^ w5551;
	assign w5596 = w5597 ^ w5579;
	assign w5638 = w5644 ^ w5596;
	assign w5640 = w5662 & w5653;
	assign w5635 = w5639 & w5638;
	assign w5708 = w47803 ^ w47801;
	assign w5709 = w47799 ^ w47797;
	assign w5710 = w47802 ^ w5708;
	assign w5786 = w47798 ^ w5710;
	assign w5783 = w47799 ^ w5710;
	assign w5711 = w47800 ^ w47798;
	assign w5715 = w47804 ^ w47798;
	assign w5785 = w5715 ^ w5710;
	assign w5797 = w47800 ^ w47797;
	assign w5792 = w5709 ^ w5715;
	assign w5789 = w5708 ^ w5797;
	assign w5788 = w47804 ^ w5789;
	assign w5725 = w47803 ^ w47802;
	assign w5790 = w5725 ^ w5792;
	assign w5793 = w5797 ^ w5725;
	assign w5799 = w47802 ^ w47800;
	assign w5784 = w5709 ^ w5799;
	assign w5795 = w47799 ^ w5715;
	assign w5791 = w47803 ^ w5795;
	assign w5685 = w47801 ^ w47802;
	assign w5671 = w5711 ^ w5709;
	assign w5787 = w5708 ^ w5671;
	assign w5670 = w5711 ^ w47799;
	assign w5794 = w47804 ^ w5670;
	assign w5798 = w47797 ^ w47803;
	assign w5796 = w47797 ^ w47802;
	assign w5782 = w5789 & w5793;
	assign w5714 = w5782 ^ w5711;
	assign w5781 = w5790 & w5788;
	assign w5780 = w5794 & w47804;
	assign w5779 = w5798 & w5783;
	assign w5713 = w5779 ^ w5709;
	assign w5778 = w5795 & w5791;
	assign w5777 = w5792 & w5785;
	assign w5776 = w5797 & w5786;
	assign w5712 = w5776 ^ w5710;
	assign w5718 = w5714 ^ w5712;
	assign w5723 = w47797 ^ w5718;
	assign w5775 = w5799 & w5784;
	assign w5732 = w5775 ^ w5781;
	assign w5773 = w5732 ^ w5723;
	assign w5684 = w5775 ^ w5776;
	assign w5731 = w5684 ^ w5685;
	assign w5730 = w5731 ^ w5713;
	assign w5772 = w5778 ^ w5730;
	assign w5774 = w5796 & w5787;
	assign w5769 = w5773 & w5772;
	assign w5842 = w47787 ^ w47785;
	assign w5843 = w47783 ^ w47781;
	assign w5844 = w47786 ^ w5842;
	assign w5920 = w47782 ^ w5844;
	assign w5917 = w47783 ^ w5844;
	assign w5845 = w47784 ^ w47782;
	assign w5849 = w47788 ^ w47782;
	assign w5919 = w5849 ^ w5844;
	assign w5931 = w47784 ^ w47781;
	assign w5926 = w5843 ^ w5849;
	assign w5923 = w5842 ^ w5931;
	assign w5922 = w47788 ^ w5923;
	assign w5859 = w47787 ^ w47786;
	assign w5924 = w5859 ^ w5926;
	assign w5927 = w5931 ^ w5859;
	assign w5933 = w47786 ^ w47784;
	assign w5918 = w5843 ^ w5933;
	assign w5929 = w47783 ^ w5849;
	assign w5925 = w47787 ^ w5929;
	assign w5819 = w47785 ^ w47786;
	assign w5805 = w5845 ^ w5843;
	assign w5921 = w5842 ^ w5805;
	assign w5804 = w5845 ^ w47783;
	assign w5928 = w47788 ^ w5804;
	assign w5932 = w47781 ^ w47787;
	assign w5930 = w47781 ^ w47786;
	assign w5916 = w5923 & w5927;
	assign w5848 = w5916 ^ w5845;
	assign w5915 = w5924 & w5922;
	assign w5914 = w5928 & w47788;
	assign w5913 = w5932 & w5917;
	assign w5847 = w5913 ^ w5843;
	assign w5912 = w5929 & w5925;
	assign w5911 = w5926 & w5919;
	assign w5910 = w5931 & w5920;
	assign w5846 = w5910 ^ w5844;
	assign w5852 = w5848 ^ w5846;
	assign w5857 = w47781 ^ w5852;
	assign w5909 = w5933 & w5918;
	assign w5866 = w5909 ^ w5915;
	assign w5907 = w5866 ^ w5857;
	assign w5818 = w5909 ^ w5910;
	assign w5865 = w5818 ^ w5819;
	assign w5864 = w5865 ^ w5847;
	assign w5906 = w5912 ^ w5864;
	assign w5908 = w5930 & w5921;
	assign w5903 = w5907 & w5906;
	assign w21423 = w47771 ^ w47769;
	assign w21424 = w47767 ^ w47765;
	assign w21425 = w47770 ^ w21423;
	assign w21501 = w47766 ^ w21425;
	assign w21498 = w47767 ^ w21425;
	assign w21426 = w47768 ^ w47766;
	assign w21430 = w47772 ^ w47766;
	assign w21500 = w21430 ^ w21425;
	assign w21512 = w47768 ^ w47765;
	assign w21507 = w21424 ^ w21430;
	assign w21504 = w21423 ^ w21512;
	assign w21503 = w47772 ^ w21504;
	assign w21440 = w47771 ^ w47770;
	assign w21505 = w21440 ^ w21507;
	assign w21508 = w21512 ^ w21440;
	assign w21514 = w47770 ^ w47768;
	assign w21499 = w21424 ^ w21514;
	assign w21510 = w47767 ^ w21430;
	assign w21506 = w47771 ^ w21510;
	assign w21400 = w47769 ^ w47770;
	assign w21386 = w21426 ^ w21424;
	assign w21502 = w21423 ^ w21386;
	assign w21385 = w21426 ^ w47767;
	assign w21509 = w47772 ^ w21385;
	assign w21513 = w47765 ^ w47771;
	assign w21511 = w47765 ^ w47770;
	assign w21497 = w21504 & w21508;
	assign w21429 = w21497 ^ w21426;
	assign w21496 = w21505 & w21503;
	assign w21495 = w21509 & w47772;
	assign w21494 = w21513 & w21498;
	assign w21428 = w21494 ^ w21424;
	assign w21493 = w21510 & w21506;
	assign w21492 = w21507 & w21500;
	assign w21491 = w21512 & w21501;
	assign w21427 = w21491 ^ w21425;
	assign w21433 = w21429 ^ w21427;
	assign w21438 = w47765 ^ w21433;
	assign w21490 = w21514 & w21499;
	assign w21447 = w21490 ^ w21496;
	assign w21488 = w21447 ^ w21438;
	assign w21399 = w21490 ^ w21491;
	assign w21446 = w21399 ^ w21400;
	assign w21445 = w21446 ^ w21428;
	assign w21487 = w21493 ^ w21445;
	assign w21489 = w21511 & w21502;
	assign w21484 = w21488 & w21487;
	assign w21557 = w47795 ^ w47793;
	assign w21558 = w47791 ^ w47789;
	assign w21559 = w47794 ^ w21557;
	assign w21635 = w47790 ^ w21559;
	assign w21632 = w47791 ^ w21559;
	assign w21560 = w47792 ^ w47790;
	assign w21564 = w47796 ^ w47790;
	assign w21634 = w21564 ^ w21559;
	assign w21646 = w47792 ^ w47789;
	assign w21641 = w21558 ^ w21564;
	assign w21638 = w21557 ^ w21646;
	assign w21637 = w47796 ^ w21638;
	assign w21574 = w47795 ^ w47794;
	assign w21639 = w21574 ^ w21641;
	assign w21642 = w21646 ^ w21574;
	assign w21648 = w47794 ^ w47792;
	assign w21633 = w21558 ^ w21648;
	assign w21644 = w47791 ^ w21564;
	assign w21640 = w47795 ^ w21644;
	assign w21534 = w47793 ^ w47794;
	assign w21520 = w21560 ^ w21558;
	assign w21636 = w21557 ^ w21520;
	assign w21519 = w21560 ^ w47791;
	assign w21643 = w47796 ^ w21519;
	assign w21647 = w47789 ^ w47795;
	assign w21645 = w47789 ^ w47794;
	assign w21631 = w21638 & w21642;
	assign w21563 = w21631 ^ w21560;
	assign w21630 = w21639 & w21637;
	assign w21629 = w21643 & w47796;
	assign w21628 = w21647 & w21632;
	assign w21562 = w21628 ^ w21558;
	assign w21627 = w21644 & w21640;
	assign w21626 = w21641 & w21634;
	assign w21625 = w21646 & w21635;
	assign w21561 = w21625 ^ w21559;
	assign w21567 = w21563 ^ w21561;
	assign w21572 = w47789 ^ w21567;
	assign w21624 = w21648 & w21633;
	assign w21581 = w21624 ^ w21630;
	assign w21622 = w21581 ^ w21572;
	assign w21533 = w21624 ^ w21625;
	assign w21580 = w21533 ^ w21534;
	assign w21579 = w21580 ^ w21562;
	assign w21621 = w21627 ^ w21579;
	assign w21623 = w21645 & w21636;
	assign w21618 = w21622 & w21621;
	assign w21691 = w47811 ^ w47809;
	assign w21692 = w47807 ^ w47805;
	assign w21693 = w47810 ^ w21691;
	assign w21769 = w47806 ^ w21693;
	assign w21766 = w47807 ^ w21693;
	assign w21694 = w47808 ^ w47806;
	assign w21698 = w47812 ^ w47806;
	assign w21768 = w21698 ^ w21693;
	assign w21780 = w47808 ^ w47805;
	assign w21775 = w21692 ^ w21698;
	assign w21772 = w21691 ^ w21780;
	assign w21771 = w47812 ^ w21772;
	assign w21708 = w47811 ^ w47810;
	assign w21773 = w21708 ^ w21775;
	assign w21776 = w21780 ^ w21708;
	assign w21782 = w47810 ^ w47808;
	assign w21767 = w21692 ^ w21782;
	assign w21778 = w47807 ^ w21698;
	assign w21774 = w47811 ^ w21778;
	assign w21668 = w47809 ^ w47810;
	assign w21654 = w21694 ^ w21692;
	assign w21770 = w21691 ^ w21654;
	assign w21653 = w21694 ^ w47807;
	assign w21777 = w47812 ^ w21653;
	assign w21781 = w47805 ^ w47811;
	assign w21779 = w47805 ^ w47810;
	assign w21765 = w21772 & w21776;
	assign w21697 = w21765 ^ w21694;
	assign w21764 = w21773 & w21771;
	assign w21763 = w21777 & w47812;
	assign w21762 = w21781 & w21766;
	assign w21696 = w21762 ^ w21692;
	assign w21761 = w21778 & w21774;
	assign w21760 = w21775 & w21768;
	assign w21759 = w21780 & w21769;
	assign w21695 = w21759 ^ w21693;
	assign w21701 = w21697 ^ w21695;
	assign w21706 = w47805 ^ w21701;
	assign w21758 = w21782 & w21767;
	assign w21715 = w21758 ^ w21764;
	assign w21756 = w21715 ^ w21706;
	assign w21667 = w21758 ^ w21759;
	assign w21714 = w21667 ^ w21668;
	assign w21713 = w21714 ^ w21696;
	assign w21755 = w21761 ^ w21713;
	assign w21757 = w21779 & w21770;
	assign w21752 = w21756 & w21755;
	assign w21825 = w47843 ^ w47841;
	assign w21826 = w47839 ^ w47837;
	assign w21827 = w47842 ^ w21825;
	assign w21903 = w47838 ^ w21827;
	assign w21900 = w47839 ^ w21827;
	assign w21828 = w47840 ^ w47838;
	assign w21832 = w47844 ^ w47838;
	assign w21902 = w21832 ^ w21827;
	assign w21914 = w47840 ^ w47837;
	assign w21909 = w21826 ^ w21832;
	assign w21906 = w21825 ^ w21914;
	assign w21905 = w47844 ^ w21906;
	assign w21842 = w47843 ^ w47842;
	assign w21907 = w21842 ^ w21909;
	assign w21910 = w21914 ^ w21842;
	assign w21916 = w47842 ^ w47840;
	assign w21901 = w21826 ^ w21916;
	assign w21912 = w47839 ^ w21832;
	assign w21908 = w47843 ^ w21912;
	assign w21802 = w47841 ^ w47842;
	assign w21788 = w21828 ^ w21826;
	assign w21904 = w21825 ^ w21788;
	assign w21787 = w21828 ^ w47839;
	assign w21911 = w47844 ^ w21787;
	assign w21915 = w47837 ^ w47843;
	assign w21913 = w47837 ^ w47842;
	assign w21899 = w21906 & w21910;
	assign w21831 = w21899 ^ w21828;
	assign w21898 = w21907 & w21905;
	assign w21897 = w21911 & w47844;
	assign w21896 = w21915 & w21900;
	assign w21830 = w21896 ^ w21826;
	assign w21895 = w21912 & w21908;
	assign w21894 = w21909 & w21902;
	assign w21893 = w21914 & w21903;
	assign w21829 = w21893 ^ w21827;
	assign w21835 = w21831 ^ w21829;
	assign w21840 = w47837 ^ w21835;
	assign w21892 = w21916 & w21901;
	assign w21849 = w21892 ^ w21898;
	assign w21890 = w21849 ^ w21840;
	assign w21801 = w21892 ^ w21893;
	assign w21848 = w21801 ^ w21802;
	assign w21847 = w21848 ^ w21830;
	assign w21889 = w21895 ^ w21847;
	assign w21891 = w21913 & w21904;
	assign w21886 = w21890 & w21889;
	assign w21959 = w47859 ^ w47857;
	assign w21960 = w47855 ^ w47853;
	assign w21961 = w47858 ^ w21959;
	assign w22037 = w47854 ^ w21961;
	assign w22034 = w47855 ^ w21961;
	assign w21962 = w47856 ^ w47854;
	assign w21966 = w47860 ^ w47854;
	assign w22036 = w21966 ^ w21961;
	assign w22048 = w47856 ^ w47853;
	assign w22043 = w21960 ^ w21966;
	assign w22040 = w21959 ^ w22048;
	assign w22039 = w47860 ^ w22040;
	assign w21976 = w47859 ^ w47858;
	assign w22041 = w21976 ^ w22043;
	assign w22044 = w22048 ^ w21976;
	assign w22050 = w47858 ^ w47856;
	assign w22035 = w21960 ^ w22050;
	assign w22046 = w47855 ^ w21966;
	assign w22042 = w47859 ^ w22046;
	assign w21936 = w47857 ^ w47858;
	assign w21922 = w21962 ^ w21960;
	assign w22038 = w21959 ^ w21922;
	assign w21921 = w21962 ^ w47855;
	assign w22045 = w47860 ^ w21921;
	assign w22049 = w47853 ^ w47859;
	assign w22047 = w47853 ^ w47858;
	assign w22033 = w22040 & w22044;
	assign w21965 = w22033 ^ w21962;
	assign w22032 = w22041 & w22039;
	assign w22031 = w22045 & w47860;
	assign w22030 = w22049 & w22034;
	assign w21964 = w22030 ^ w21960;
	assign w22029 = w22046 & w22042;
	assign w22028 = w22043 & w22036;
	assign w22027 = w22048 & w22037;
	assign w21963 = w22027 ^ w21961;
	assign w21969 = w21965 ^ w21963;
	assign w21974 = w47853 ^ w21969;
	assign w22026 = w22050 & w22035;
	assign w21983 = w22026 ^ w22032;
	assign w22024 = w21983 ^ w21974;
	assign w21935 = w22026 ^ w22027;
	assign w21982 = w21935 ^ w21936;
	assign w21981 = w21982 ^ w21964;
	assign w22023 = w22029 ^ w21981;
	assign w22025 = w22047 & w22038;
	assign w22020 = w22024 & w22023;
	assign w25845 = w47827 ^ w47825;
	assign w25846 = w47823 ^ w47821;
	assign w25847 = w47826 ^ w25845;
	assign w25923 = w47822 ^ w25847;
	assign w25920 = w47823 ^ w25847;
	assign w25848 = w47824 ^ w47822;
	assign w25852 = w47828 ^ w47822;
	assign w25922 = w25852 ^ w25847;
	assign w25934 = w47824 ^ w47821;
	assign w25929 = w25846 ^ w25852;
	assign w25926 = w25845 ^ w25934;
	assign w25925 = w47828 ^ w25926;
	assign w25862 = w47827 ^ w47826;
	assign w25927 = w25862 ^ w25929;
	assign w25930 = w25934 ^ w25862;
	assign w25936 = w47826 ^ w47824;
	assign w25921 = w25846 ^ w25936;
	assign w25932 = w47823 ^ w25852;
	assign w25928 = w47827 ^ w25932;
	assign w25822 = w47825 ^ w47826;
	assign w25808 = w25848 ^ w25846;
	assign w25924 = w25845 ^ w25808;
	assign w25807 = w25848 ^ w47823;
	assign w25931 = w47828 ^ w25807;
	assign w25935 = w47821 ^ w47827;
	assign w25933 = w47821 ^ w47826;
	assign w25919 = w25926 & w25930;
	assign w25851 = w25919 ^ w25848;
	assign w25918 = w25927 & w25925;
	assign w25917 = w25931 & w47828;
	assign w25916 = w25935 & w25920;
	assign w25850 = w25916 ^ w25846;
	assign w25915 = w25932 & w25928;
	assign w25914 = w25929 & w25922;
	assign w25913 = w25934 & w25923;
	assign w25849 = w25913 ^ w25847;
	assign w25855 = w25851 ^ w25849;
	assign w25860 = w47821 ^ w25855;
	assign w25912 = w25936 & w25921;
	assign w25869 = w25912 ^ w25918;
	assign w25910 = w25869 ^ w25860;
	assign w25821 = w25912 ^ w25913;
	assign w25868 = w25821 ^ w25822;
	assign w25867 = w25868 ^ w25850;
	assign w25909 = w25915 ^ w25867;
	assign w25911 = w25933 & w25924;
	assign w25906 = w25910 & w25909;
	assign w28927 = w47779 ^ w47777;
	assign w28928 = w47775 ^ w47773;
	assign w28929 = w47778 ^ w28927;
	assign w29005 = w47774 ^ w28929;
	assign w29002 = w47775 ^ w28929;
	assign w28930 = w47776 ^ w47774;
	assign w28934 = w47780 ^ w47774;
	assign w29004 = w28934 ^ w28929;
	assign w29016 = w47776 ^ w47773;
	assign w29011 = w28928 ^ w28934;
	assign w29008 = w28927 ^ w29016;
	assign w29007 = w47780 ^ w29008;
	assign w28944 = w47779 ^ w47778;
	assign w29009 = w28944 ^ w29011;
	assign w29012 = w29016 ^ w28944;
	assign w29018 = w47778 ^ w47776;
	assign w29003 = w28928 ^ w29018;
	assign w29014 = w47775 ^ w28934;
	assign w29010 = w47779 ^ w29014;
	assign w28904 = w47777 ^ w47778;
	assign w28890 = w28930 ^ w28928;
	assign w29006 = w28927 ^ w28890;
	assign w28889 = w28930 ^ w47775;
	assign w29013 = w47780 ^ w28889;
	assign w29017 = w47773 ^ w47779;
	assign w29015 = w47773 ^ w47778;
	assign w29001 = w29008 & w29012;
	assign w28933 = w29001 ^ w28930;
	assign w29000 = w29009 & w29007;
	assign w28999 = w29013 & w47780;
	assign w28998 = w29017 & w29002;
	assign w28932 = w28998 ^ w28928;
	assign w28997 = w29014 & w29010;
	assign w28996 = w29011 & w29004;
	assign w28995 = w29016 & w29005;
	assign w28931 = w28995 ^ w28929;
	assign w28937 = w28933 ^ w28931;
	assign w28942 = w47773 ^ w28937;
	assign w28994 = w29018 & w29003;
	assign w28951 = w28994 ^ w29000;
	assign w28992 = w28951 ^ w28942;
	assign w28903 = w28994 ^ w28995;
	assign w28950 = w28903 ^ w28904;
	assign w28949 = w28950 ^ w28932;
	assign w28991 = w28997 ^ w28949;
	assign w28993 = w29015 & w29006;
	assign w28988 = w28992 & w28991;
	assign w32545 = w47835 ^ w47833;
	assign w32546 = w47831 ^ w47829;
	assign w32547 = w47834 ^ w32545;
	assign w32623 = w47830 ^ w32547;
	assign w32620 = w47831 ^ w32547;
	assign w32548 = w47832 ^ w47830;
	assign w32552 = w47836 ^ w47830;
	assign w32622 = w32552 ^ w32547;
	assign w32634 = w47832 ^ w47829;
	assign w32629 = w32546 ^ w32552;
	assign w32626 = w32545 ^ w32634;
	assign w32625 = w47836 ^ w32626;
	assign w32562 = w47835 ^ w47834;
	assign w32627 = w32562 ^ w32629;
	assign w32630 = w32634 ^ w32562;
	assign w32636 = w47834 ^ w47832;
	assign w32621 = w32546 ^ w32636;
	assign w32632 = w47831 ^ w32552;
	assign w32628 = w47835 ^ w32632;
	assign w32522 = w47833 ^ w47834;
	assign w32508 = w32548 ^ w32546;
	assign w32624 = w32545 ^ w32508;
	assign w32507 = w32548 ^ w47831;
	assign w32631 = w47836 ^ w32507;
	assign w32635 = w47829 ^ w47835;
	assign w32633 = w47829 ^ w47834;
	assign w32619 = w32626 & w32630;
	assign w32551 = w32619 ^ w32548;
	assign w32618 = w32627 & w32625;
	assign w32617 = w32631 & w47836;
	assign w32616 = w32635 & w32620;
	assign w32550 = w32616 ^ w32546;
	assign w32615 = w32632 & w32628;
	assign w32614 = w32629 & w32622;
	assign w32613 = w32634 & w32623;
	assign w32549 = w32613 ^ w32547;
	assign w32555 = w32551 ^ w32549;
	assign w32560 = w47829 ^ w32555;
	assign w32612 = w32636 & w32621;
	assign w32569 = w32612 ^ w32618;
	assign w32610 = w32569 ^ w32560;
	assign w32521 = w32612 ^ w32613;
	assign w32568 = w32521 ^ w32522;
	assign w32567 = w32568 ^ w32550;
	assign w32609 = w32615 ^ w32567;
	assign w32611 = w32633 & w32624;
	assign w32606 = w32610 & w32609;
	assign w36029 = w47819 ^ w47817;
	assign w36030 = w47815 ^ w47813;
	assign w36031 = w47818 ^ w36029;
	assign w36107 = w47814 ^ w36031;
	assign w36104 = w47815 ^ w36031;
	assign w36032 = w47816 ^ w47814;
	assign w36036 = w47820 ^ w47814;
	assign w36106 = w36036 ^ w36031;
	assign w36118 = w47816 ^ w47813;
	assign w36113 = w36030 ^ w36036;
	assign w36110 = w36029 ^ w36118;
	assign w36109 = w47820 ^ w36110;
	assign w36046 = w47819 ^ w47818;
	assign w36111 = w36046 ^ w36113;
	assign w36114 = w36118 ^ w36046;
	assign w36120 = w47818 ^ w47816;
	assign w36105 = w36030 ^ w36120;
	assign w36116 = w47815 ^ w36036;
	assign w36112 = w47819 ^ w36116;
	assign w36006 = w47817 ^ w47818;
	assign w35992 = w36032 ^ w36030;
	assign w36108 = w36029 ^ w35992;
	assign w35991 = w36032 ^ w47815;
	assign w36115 = w47820 ^ w35991;
	assign w36119 = w47813 ^ w47819;
	assign w36117 = w47813 ^ w47818;
	assign w36103 = w36110 & w36114;
	assign w36035 = w36103 ^ w36032;
	assign w36102 = w36111 & w36109;
	assign w36101 = w36115 & w47820;
	assign w36100 = w36119 & w36104;
	assign w36034 = w36100 ^ w36030;
	assign w36099 = w36116 & w36112;
	assign w36098 = w36113 & w36106;
	assign w36097 = w36118 & w36107;
	assign w36033 = w36097 ^ w36031;
	assign w36039 = w36035 ^ w36033;
	assign w36044 = w47813 ^ w36039;
	assign w36096 = w36120 & w36105;
	assign w36053 = w36096 ^ w36102;
	assign w36094 = w36053 ^ w36044;
	assign w36005 = w36096 ^ w36097;
	assign w36052 = w36005 ^ w36006;
	assign w36051 = w36052 ^ w36034;
	assign w36093 = w36099 ^ w36051;
	assign w36095 = w36117 & w36108;
	assign w36090 = w36094 & w36093;
	assign w38575 = w47891 ^ w47889;
	assign w38576 = w47887 ^ w47885;
	assign w38577 = w47890 ^ w38575;
	assign w38653 = w47886 ^ w38577;
	assign w38650 = w47887 ^ w38577;
	assign w38578 = w47888 ^ w47886;
	assign w38582 = w47892 ^ w47886;
	assign w38652 = w38582 ^ w38577;
	assign w38664 = w47888 ^ w47885;
	assign w38659 = w38576 ^ w38582;
	assign w38656 = w38575 ^ w38664;
	assign w38655 = w47892 ^ w38656;
	assign w38592 = w47891 ^ w47890;
	assign w38657 = w38592 ^ w38659;
	assign w38660 = w38664 ^ w38592;
	assign w38666 = w47890 ^ w47888;
	assign w38651 = w38576 ^ w38666;
	assign w38662 = w47887 ^ w38582;
	assign w38658 = w47891 ^ w38662;
	assign w38552 = w47889 ^ w47890;
	assign w38538 = w38578 ^ w38576;
	assign w38654 = w38575 ^ w38538;
	assign w38537 = w38578 ^ w47887;
	assign w38661 = w47892 ^ w38537;
	assign w38665 = w47885 ^ w47891;
	assign w38663 = w47885 ^ w47890;
	assign w38649 = w38656 & w38660;
	assign w38581 = w38649 ^ w38578;
	assign w38648 = w38657 & w38655;
	assign w38647 = w38661 & w47892;
	assign w38646 = w38665 & w38650;
	assign w38580 = w38646 ^ w38576;
	assign w38645 = w38662 & w38658;
	assign w38644 = w38659 & w38652;
	assign w38643 = w38664 & w38653;
	assign w38579 = w38643 ^ w38577;
	assign w38585 = w38581 ^ w38579;
	assign w38590 = w47885 ^ w38585;
	assign w38642 = w38666 & w38651;
	assign w38599 = w38642 ^ w38648;
	assign w38640 = w38599 ^ w38590;
	assign w38551 = w38642 ^ w38643;
	assign w38598 = w38551 ^ w38552;
	assign w38597 = w38598 ^ w38580;
	assign w38639 = w38645 ^ w38597;
	assign w38641 = w38663 & w38654;
	assign w38636 = w38640 & w38639;
	assign w43682 = w3627 ^ w3633;
	assign w3530 = w43682 ^ w3546;
	assign w3623 = w3536 ^ w3530;
	assign w3569 = w3537 ^ w43682;
	assign w3525 = w21 ^ w3569;
	assign w3617 = w3622 ^ w3525;
	assign w43683 = w3627 ^ w3630;
	assign w3527 = w3628 ^ w43683;
	assign w3572 = w3631 ^ w3527;
	assign w3618 = w17 ^ w3572;
	assign w3616 = w3617 & w3618;
	assign w3614 = w3622 ^ w3616;
	assign w3573 = w3616 ^ w3527;
	assign w3574 = w3616 ^ w3633;
	assign w3579 = w3574 ^ w3630;
	assign w3568 = w3542 ^ w43683;
	assign w3624 = w3568 ^ w3543;
	assign w3615 = w3616 ^ w3624;
	assign w3621 = w3622 ^ w3624;
	assign w3620 = w3623 & w3621;
	assign w3619 = w3620 ^ w3525;
	assign w3577 = w3620 ^ w3632;
	assign w3581 = w3577 ^ w3541;
	assign w3578 = w23 ^ w3581;
	assign w3607 = w3579 ^ w3578;
	assign w3580 = w3620 ^ w3531;
	assign w3582 = w21 ^ w3581;
	assign w3613 = w3624 & w3614;
	assign w3611 = w3613 ^ w3621;
	assign w3610 = w3619 & w3611;
	assign w3532 = w3610 ^ w3536;
	assign w3609 = w3532 ^ w3530;
	assign w3575 = w3610 ^ w3634;
	assign w3606 = w3532 ^ w3580;
	assign w3601 = w3615 & w16;
	assign w3600 = w3606 & w3636;
	assign w3599 = w3609 & w3648;
	assign w3598 = w3619 & w3638;
	assign w3566 = w3598 ^ w3599;
	assign w3597 = w3607 & w3639;
	assign w3592 = w3615 & w3647;
	assign w3591 = w3606 & w3651;
	assign w3550 = w3600 ^ w3591;
	assign w3590 = w3609 & w3644;
	assign w3548 = w3598 ^ w3590;
	assign w3589 = w3619 & w3645;
	assign w3588 = w3607 & w3650;
	assign w43684 = w3599 ^ w3600;
	assign w43686 = w3613 ^ w3631;
	assign w3605 = w43686 ^ w3524;
	assign w3603 = w3605 & w3642;
	assign w3594 = w3605 & w3646;
	assign w43685 = w3601 ^ w3603;
	assign w3535 = w17 ^ w43686;
	assign w3612 = w3535 ^ w3573;
	assign w3583 = w3535 ^ w3575;
	assign w3576 = w3546 ^ w3583;
	assign w3608 = w3579 ^ w3576;
	assign w3604 = w3583 ^ w3582;
	assign w3602 = w3612 & w3641;
	assign w3596 = w3604 & w3637;
	assign w3526 = w3596 ^ w43684;
	assign w3551 = w3596 ^ w3599;
	assign w3554 = ~w3551;
	assign w3555 = w3596 ^ w3597;
	assign w3561 = w3592 ^ w3526;
	assign w3564 = ~w3561;
	assign w3567 = w3597 ^ w3526;
	assign w3595 = w3608 & w3640;
	assign w3534 = w3591 ^ w3595;
	assign w3557 = ~w3534;
	assign w3558 = w3557 ^ w3589;
	assign w3562 = w3558 ^ w43685;
	assign w3559 = w3588 ^ w3562;
	assign w3593 = w3612 & w3643;
	assign w3587 = w3604 & w3652;
	assign w3586 = w3608 & w3649;
	assign w3556 = w3597 ^ w3586;
	assign w3560 = ~w3556;
	assign w3653 = w3560 ^ w3559;
	assign w47922 = ~w3653;
	assign w1911 = w253 ^ w47922;
	assign w1943 = w221 ^ w1911;
	assign w1975 = w189 ^ w1943;
	assign w2007 = w157 ^ w1975;
	assign w43516 = w3587 ^ w3588;
	assign w3552 = w3548 ^ w43516;
	assign w3549 = w43685 ^ w3552;
	assign w3656 = w3550 ^ w3549;
	assign w3553 = w3557 ^ w3552;
	assign w3655 = w3554 ^ w3553;
	assign w47917 = ~w3656;
	assign w47918 = ~w3655;
	assign w1907 = w249 ^ w47918;
	assign w1939 = w217 ^ w1907;
	assign w2042 = w248 ^ w47917;
	assign w1971 = w185 ^ w1939;
	assign w2003 = w153 ^ w1971;
	assign w3539 = w3593 ^ w43516;
	assign w3538 = w3594 ^ w3539;
	assign w3533 = w3602 ^ w3538;
	assign w3528 = w3603 ^ w3533;
	assign w47921 = w43684 ^ w3528;
	assign w3654 = w3528 ^ w3555;
	assign w3563 = w3539 ^ w3562;
	assign w47919 = w3564 ^ w3563;
	assign w3565 = w3601 ^ w3533;
	assign w47920 = w3566 ^ w3565;
	assign w47924 = w3538 ^ w3567;
	assign w47923 = ~w3654;
	assign w1912 = w254 ^ w47923;
	assign w1910 = w252 ^ w47921;
	assign w1909 = w251 ^ w47920;
	assign w1941 = w219 ^ w1909;
	assign w1913 = w255 ^ w47924;
	assign w1945 = w223 ^ w1913;
	assign w1908 = w250 ^ w47919;
	assign w1942 = w220 ^ w1910;
	assign w1944 = w222 ^ w1912;
	assign w1940 = w218 ^ w1908;
	assign w1976 = w190 ^ w1944;
	assign w2008 = w158 ^ w1976;
	assign w1977 = w191 ^ w1945;
	assign w2009 = w159 ^ w1977;
	assign w1974 = w188 ^ w1942;
	assign w2006 = w156 ^ w1974;
	assign w1973 = w187 ^ w1941;
	assign w2005 = w155 ^ w1973;
	assign w1972 = w186 ^ w1940;
	assign w2004 = w154 ^ w1972;
	assign w4097 = w2003 ^ w2005;
	assign w4098 = w2007 ^ w2009;
	assign w4099 = w2004 ^ w4097;
	assign w4176 = w2008 ^ w4099;
	assign w4173 = w2007 ^ w4099;
	assign w4100 = w2006 ^ w2008;
	assign w4187 = w2006 ^ w2009;
	assign w4179 = w4097 ^ w4187;
	assign w4114 = w2003 ^ w2004;
	assign w4183 = w4187 ^ w4114;
	assign w4189 = w2004 ^ w2006;
	assign w4174 = w4098 ^ w4189;
	assign w4074 = w2005 ^ w2004;
	assign w4060 = w4100 ^ w4098;
	assign w4177 = w4097 ^ w4060;
	assign w4059 = w4100 ^ w2007;
	assign w4188 = w2009 ^ w2003;
	assign w4186 = w2009 ^ w2004;
	assign w4172 = w4179 & w4183;
	assign w4103 = w4172 ^ w4100;
	assign w4169 = w4188 & w4173;
	assign w4102 = w4169 ^ w4098;
	assign w4166 = w4187 & w4176;
	assign w4101 = w4166 ^ w4099;
	assign w4107 = w4103 ^ w4101;
	assign w4112 = w2009 ^ w4107;
	assign w4165 = w4189 & w4174;
	assign w4073 = w4165 ^ w4166;
	assign w4120 = w4073 ^ w4074;
	assign w4119 = w4120 ^ w4102;
	assign w4164 = w4186 & w4177;
	assign w43687 = w3761 ^ w3767;
	assign w3673 = w3705 ^ w43687;
	assign w3716 = w13 ^ w3673;
	assign w3751 = w3756 ^ w3716;
	assign w3711 = w43687 ^ w3696;
	assign w3757 = w3719 ^ w3711;
	assign w43688 = w3761 ^ w3764;
	assign w3714 = w3762 ^ w43688;
	assign w3670 = w3765 ^ w3714;
	assign w3752 = w9 ^ w3670;
	assign w3750 = w3751 & w3752;
	assign w3748 = w3756 ^ w3750;
	assign w3669 = w3750 ^ w3714;
	assign w3668 = w3750 ^ w3767;
	assign w3663 = w3668 ^ w3764;
	assign w3674 = w3700 ^ w43688;
	assign w3758 = w3674 ^ w3699;
	assign w3749 = w3750 ^ w3758;
	assign w3755 = w3756 ^ w3758;
	assign w3754 = w3757 & w3755;
	assign w3753 = w3754 ^ w3716;
	assign w3665 = w3754 ^ w3766;
	assign w3661 = w3665 ^ w3701;
	assign w3664 = w15 ^ w3661;
	assign w3741 = w3663 ^ w3664;
	assign w3662 = w3754 ^ w3710;
	assign w3660 = w13 ^ w3661;
	assign w3747 = w3758 & w3748;
	assign w3745 = w3747 ^ w3755;
	assign w3744 = w3753 & w3745;
	assign w3709 = w3744 ^ w3719;
	assign w3743 = w3709 ^ w3711;
	assign w3667 = w3744 ^ w3768;
	assign w3740 = w3709 ^ w3662;
	assign w3735 = w3749 & w8;
	assign w3734 = w3740 & w3770;
	assign w3733 = w3743 & w3782;
	assign w3732 = w3753 & w3772;
	assign w3676 = w3732 ^ w3733;
	assign w3731 = w3741 & w3773;
	assign w3726 = w3749 & w3781;
	assign w3725 = w3740 & w3785;
	assign w3692 = w3734 ^ w3725;
	assign w3724 = w3743 & w3778;
	assign w3694 = w3732 ^ w3724;
	assign w3723 = w3753 & w3779;
	assign w3722 = w3741 & w3784;
	assign w43690 = w3733 ^ w3734;
	assign w43692 = w3747 ^ w3765;
	assign w3739 = w43692 ^ w3717;
	assign w3737 = w3739 & w3776;
	assign w3728 = w3739 & w3780;
	assign w43691 = w3735 ^ w3737;
	assign w3706 = w9 ^ w43692;
	assign w3746 = w3706 ^ w3669;
	assign w3659 = w3706 ^ w3667;
	assign w3666 = w3696 ^ w3659;
	assign w3742 = w3663 ^ w3666;
	assign w3738 = w3659 ^ w3660;
	assign w3736 = w3746 & w3775;
	assign w3730 = w3738 & w3771;
	assign w3715 = w3730 ^ w43690;
	assign w3691 = w3730 ^ w3733;
	assign w3688 = ~w3691;
	assign w3687 = w3730 ^ w3731;
	assign w3681 = w3726 ^ w3715;
	assign w3678 = ~w3681;
	assign w3675 = w3731 ^ w3715;
	assign w3729 = w3742 & w3774;
	assign w3707 = w3725 ^ w3729;
	assign w3685 = ~w3707;
	assign w3684 = w3685 ^ w3723;
	assign w3680 = w3684 ^ w43691;
	assign w3683 = w3722 ^ w3680;
	assign w3727 = w3746 & w3777;
	assign w3721 = w3738 & w3786;
	assign w3720 = w3742 & w3783;
	assign w3686 = w3731 ^ w3720;
	assign w3682 = ~w3686;
	assign w3787 = w3682 ^ w3683;
	assign w47914 = ~w3787;
	assign w1904 = w245 ^ w47914;
	assign w1935 = w213 ^ w1904;
	assign w1967 = w181 ^ w1935;
	assign w1999 = w149 ^ w1967;
	assign w43689 = w3721 ^ w3722;
	assign w3703 = w3727 ^ w43689;
	assign w3704 = w3728 ^ w3703;
	assign w3708 = w3736 ^ w3704;
	assign w3713 = w3737 ^ w3708;
	assign w47913 = w43690 ^ w3713;
	assign w3788 = w3713 ^ w3687;
	assign w3679 = w3703 ^ w3680;
	assign w47911 = w3678 ^ w3679;
	assign w3677 = w3735 ^ w3708;
	assign w47912 = w3676 ^ w3677;
	assign w47916 = w3704 ^ w3675;
	assign w47915 = ~w3788;
	assign w1906 = w247 ^ w47916;
	assign w1937 = w215 ^ w1906;
	assign w1905 = w246 ^ w47915;
	assign w1936 = w214 ^ w1905;
	assign w1903 = w244 ^ w47913;
	assign w1934 = w212 ^ w1903;
	assign w1902 = w243 ^ w47912;
	assign w1901 = w242 ^ w47911;
	assign w1932 = w210 ^ w1901;
	assign w1933 = w211 ^ w1902;
	assign w1969 = w183 ^ w1937;
	assign w1968 = w182 ^ w1936;
	assign w1966 = w180 ^ w1934;
	assign w1965 = w179 ^ w1933;
	assign w1964 = w178 ^ w1932;
	assign w1998 = w148 ^ w1966;
	assign w2001 = w151 ^ w1969;
	assign w4233 = w1999 ^ w2001;
	assign w4321 = w1998 ^ w2001;
	assign w2000 = w150 ^ w1968;
	assign w4235 = w1998 ^ w2000;
	assign w4195 = w4235 ^ w4233;
	assign w4194 = w4235 ^ w1999;
	assign w1997 = w147 ^ w1965;
	assign w1996 = w146 ^ w1964;
	assign w4323 = w1996 ^ w1998;
	assign w4308 = w4233 ^ w4323;
	assign w4209 = w1997 ^ w1996;
	assign w4320 = w2001 ^ w1996;
	assign w4299 = w4323 & w4308;
	assign w3690 = w3694 ^ w43689;
	assign w3693 = w43691 ^ w3690;
	assign w3790 = w3692 ^ w3693;
	assign w3689 = w3685 ^ w3690;
	assign w3789 = w3688 ^ w3689;
	assign w47909 = ~w3790;
	assign w47910 = ~w3789;
	assign w1900 = w241 ^ w47910;
	assign w1931 = w209 ^ w1900;
	assign w1899 = w240 ^ w47909;
	assign w1930 = w208 ^ w1899;
	assign w1963 = w177 ^ w1931;
	assign w1962 = w176 ^ w1930;
	assign w1995 = w145 ^ w1963;
	assign w4232 = w1995 ^ w1997;
	assign w4234 = w1996 ^ w4232;
	assign w4310 = w2000 ^ w4234;
	assign w4307 = w1999 ^ w4234;
	assign w4313 = w4232 ^ w4321;
	assign w4249 = w1995 ^ w1996;
	assign w4317 = w4321 ^ w4249;
	assign w4311 = w4232 ^ w4195;
	assign w4322 = w2001 ^ w1995;
	assign w4306 = w4313 & w4317;
	assign w4238 = w4306 ^ w4235;
	assign w4303 = w4322 & w4307;
	assign w4237 = w4303 ^ w4233;
	assign w4300 = w4321 & w4310;
	assign w4236 = w4300 ^ w4234;
	assign w4242 = w4238 ^ w4236;
	assign w4247 = w2001 ^ w4242;
	assign w4208 = w4299 ^ w4300;
	assign w4255 = w4208 ^ w4209;
	assign w4254 = w4255 ^ w4237;
	assign w4298 = w4320 & w4311;
	assign w1994 = w144 ^ w1962;
	assign w4312 = w1994 ^ w4313;
	assign w4239 = w1994 ^ w2000;
	assign w4309 = w4239 ^ w4234;
	assign w4316 = w4233 ^ w4239;
	assign w4314 = w4249 ^ w4316;
	assign w4319 = w1999 ^ w4239;
	assign w4315 = w1995 ^ w4319;
	assign w4318 = w1994 ^ w4194;
	assign w4305 = w4314 & w4312;
	assign w4256 = w4299 ^ w4305;
	assign w4297 = w4256 ^ w4247;
	assign w4304 = w4318 & w1994;
	assign w4302 = w4319 & w4315;
	assign w4296 = w4302 ^ w4254;
	assign w4301 = w4316 & w4309;
	assign w4293 = w4297 & w4296;
	assign w43693 = w3895 ^ w3898;
	assign w3808 = w3834 ^ w43693;
	assign w3892 = w3808 ^ w3833;
	assign w3889 = w3890 ^ w3892;
	assign w3848 = w3896 ^ w43693;
	assign w3804 = w3899 ^ w3848;
	assign w3886 = w1 ^ w3804;
	assign w43696 = w3895 ^ w3901;
	assign w3807 = w3839 ^ w43696;
	assign w3850 = w5 ^ w3807;
	assign w3885 = w3890 ^ w3850;
	assign w3884 = w3885 & w3886;
	assign w3883 = w3884 ^ w3892;
	assign w3882 = w3890 ^ w3884;
	assign w3803 = w3884 ^ w3848;
	assign w3802 = w3884 ^ w3901;
	assign w3797 = w3802 ^ w3898;
	assign w3881 = w3892 & w3882;
	assign w3879 = w3881 ^ w3889;
	assign w3869 = w3883 & w0;
	assign w3860 = w3883 & w3915;
	assign w43695 = w3881 ^ w3899;
	assign w3873 = w43695 ^ w3851;
	assign w3871 = w3873 & w3910;
	assign w3862 = w3873 & w3914;
	assign w3840 = w1 ^ w43695;
	assign w3880 = w3840 ^ w3803;
	assign w3870 = w3880 & w3909;
	assign w3861 = w3880 & w3911;
	assign w3845 = w43696 ^ w3830;
	assign w3891 = w3853 ^ w3845;
	assign w3888 = w3891 & w3889;
	assign w3887 = w3888 ^ w3850;
	assign w3799 = w3888 ^ w3900;
	assign w3795 = w3799 ^ w3835;
	assign w3798 = w7 ^ w3795;
	assign w3875 = w3797 ^ w3798;
	assign w3796 = w3888 ^ w3844;
	assign w3794 = w5 ^ w3795;
	assign w3878 = w3887 & w3879;
	assign w3843 = w3878 ^ w3853;
	assign w3877 = w3843 ^ w3845;
	assign w3801 = w3878 ^ w3902;
	assign w3793 = w3840 ^ w3801;
	assign w3800 = w3830 ^ w3793;
	assign w3876 = w3797 ^ w3800;
	assign w3874 = w3843 ^ w3796;
	assign w3872 = w3793 ^ w3794;
	assign w3868 = w3874 & w3904;
	assign w3867 = w3877 & w3916;
	assign w3866 = w3887 & w3906;
	assign w3810 = w3866 ^ w3867;
	assign w3865 = w3875 & w3907;
	assign w3864 = w3872 & w3905;
	assign w3825 = w3864 ^ w3867;
	assign w3822 = ~w3825;
	assign w3821 = w3864 ^ w3865;
	assign w3863 = w3876 & w3908;
	assign w3859 = w3874 & w3919;
	assign w3841 = w3859 ^ w3863;
	assign w3826 = w3868 ^ w3859;
	assign w3819 = ~w3841;
	assign w3858 = w3877 & w3912;
	assign w3828 = w3866 ^ w3858;
	assign w3857 = w3887 & w3913;
	assign w3818 = w3819 ^ w3857;
	assign w3856 = w3875 & w3918;
	assign w3855 = w3872 & w3920;
	assign w3854 = w3876 & w3917;
	assign w3820 = w3865 ^ w3854;
	assign w3816 = ~w3820;
	assign w43694 = w3855 ^ w3856;
	assign w3837 = w3861 ^ w43694;
	assign w3838 = w3862 ^ w3837;
	assign w3842 = w3870 ^ w3838;
	assign w3847 = w3871 ^ w3842;
	assign w3922 = w3847 ^ w3821;
	assign w3811 = w3869 ^ w3842;
	assign w47904 = w3810 ^ w3811;
	assign w1894 = w235 ^ w47904;
	assign w47907 = ~w3922;
	assign w1897 = w238 ^ w47907;
	assign w1928 = w206 ^ w1897;
	assign w1925 = w203 ^ w1894;
	assign w1957 = w171 ^ w1925;
	assign w1960 = w174 ^ w1928;
	assign w1989 = w139 ^ w1957;
	assign w1992 = w142 ^ w1960;
	assign w3824 = w3828 ^ w43694;
	assign w3823 = w3819 ^ w3824;
	assign w3923 = w3822 ^ w3823;
	assign w47902 = ~w3923;
	assign w1892 = w233 ^ w47902;
	assign w1923 = w201 ^ w1892;
	assign w1955 = w169 ^ w1923;
	assign w1987 = w137 ^ w1955;
	assign w4366 = w1987 ^ w1989;
	assign w43697 = w3867 ^ w3868;
	assign w47905 = w43697 ^ w3847;
	assign w1895 = w236 ^ w47905;
	assign w1926 = w204 ^ w1895;
	assign w1958 = w172 ^ w1926;
	assign w1990 = w140 ^ w1958;
	assign w4369 = w1990 ^ w1992;
	assign w3849 = w3864 ^ w43697;
	assign w3815 = w3860 ^ w3849;
	assign w3812 = ~w3815;
	assign w3809 = w3865 ^ w3849;
	assign w47908 = w3838 ^ w3809;
	assign w1898 = w239 ^ w47908;
	assign w1929 = w207 ^ w1898;
	assign w1961 = w175 ^ w1929;
	assign w1993 = w143 ^ w1961;
	assign w4455 = w1990 ^ w1993;
	assign w4447 = w4366 ^ w4455;
	assign w4456 = w1993 ^ w1987;
	assign w43698 = w3869 ^ w3871;
	assign w3827 = w43698 ^ w3824;
	assign w3924 = w3826 ^ w3827;
	assign w47901 = ~w3924;
	assign w1891 = w232 ^ w47901;
	assign w1922 = w200 ^ w1891;
	assign w1954 = w168 ^ w1922;
	assign w1986 = w136 ^ w1954;
	assign w4373 = w1986 ^ w1992;
	assign w4446 = w1986 ^ w4447;
	assign w3814 = w3818 ^ w43698;
	assign w3817 = w3856 ^ w3814;
	assign w3921 = w3816 ^ w3817;
	assign w3813 = w3837 ^ w3814;
	assign w47903 = w3812 ^ w3813;
	assign w1893 = w234 ^ w47903;
	assign w47906 = ~w3921;
	assign w1896 = w237 ^ w47906;
	assign w1927 = w205 ^ w1896;
	assign w1959 = w173 ^ w1927;
	assign w1924 = w202 ^ w1893;
	assign w1956 = w170 ^ w1924;
	assign w1991 = w141 ^ w1959;
	assign w4367 = w1991 ^ w1993;
	assign w4450 = w4367 ^ w4373;
	assign w4453 = w1991 ^ w4373;
	assign w4449 = w1987 ^ w4453;
	assign w4329 = w4369 ^ w4367;
	assign w4445 = w4366 ^ w4329;
	assign w4328 = w4369 ^ w1991;
	assign w4452 = w1986 ^ w4328;
	assign w4438 = w4452 & w1986;
	assign w4436 = w4453 & w4449;
	assign w1988 = w138 ^ w1956;
	assign w4368 = w1988 ^ w4366;
	assign w4444 = w1992 ^ w4368;
	assign w4441 = w1991 ^ w4368;
	assign w4443 = w4373 ^ w4368;
	assign w4383 = w1987 ^ w1988;
	assign w4448 = w4383 ^ w4450;
	assign w4451 = w4455 ^ w4383;
	assign w4457 = w1988 ^ w1990;
	assign w4442 = w4367 ^ w4457;
	assign w4343 = w1989 ^ w1988;
	assign w4454 = w1993 ^ w1988;
	assign w4440 = w4447 & w4451;
	assign w4372 = w4440 ^ w4369;
	assign w4439 = w4448 & w4446;
	assign w4437 = w4456 & w4441;
	assign w4371 = w4437 ^ w4367;
	assign w4435 = w4450 & w4443;
	assign w4434 = w4455 & w4444;
	assign w4370 = w4434 ^ w4368;
	assign w4376 = w4372 ^ w4370;
	assign w4381 = w1993 ^ w4376;
	assign w4433 = w4457 & w4442;
	assign w4390 = w4433 ^ w4439;
	assign w4431 = w4390 ^ w4381;
	assign w4342 = w4433 ^ w4434;
	assign w4389 = w4342 ^ w4343;
	assign w4388 = w4389 ^ w4371;
	assign w4430 = w4436 ^ w4388;
	assign w4432 = w4454 & w4445;
	assign w4427 = w4431 & w4430;
	assign w43699 = w4029 ^ w4035;
	assign w3979 = w43699 ^ w3964;
	assign w4025 = w3987 ^ w3979;
	assign w3941 = w3973 ^ w43699;
	assign w3984 = w29 ^ w3941;
	assign w4019 = w4024 ^ w3984;
	assign w43700 = w4029 ^ w4032;
	assign w3982 = w4030 ^ w43700;
	assign w3938 = w4033 ^ w3982;
	assign w4020 = w25 ^ w3938;
	assign w4018 = w4019 & w4020;
	assign w4016 = w4024 ^ w4018;
	assign w3937 = w4018 ^ w3982;
	assign w3936 = w4018 ^ w4035;
	assign w3931 = w3936 ^ w4032;
	assign w3942 = w3968 ^ w43700;
	assign w4026 = w3942 ^ w3967;
	assign w4017 = w4018 ^ w4026;
	assign w4023 = w4024 ^ w4026;
	assign w4022 = w4025 & w4023;
	assign w4021 = w4022 ^ w3984;
	assign w3933 = w4022 ^ w4034;
	assign w3929 = w3933 ^ w3969;
	assign w3932 = w31 ^ w3929;
	assign w4009 = w3931 ^ w3932;
	assign w3930 = w4022 ^ w3978;
	assign w3928 = w29 ^ w3929;
	assign w4015 = w4026 & w4016;
	assign w4013 = w4015 ^ w4023;
	assign w4012 = w4021 & w4013;
	assign w3977 = w4012 ^ w3987;
	assign w4011 = w3977 ^ w3979;
	assign w3935 = w4012 ^ w4036;
	assign w4008 = w3977 ^ w3930;
	assign w4003 = w4017 & w24;
	assign w4002 = w4008 & w4038;
	assign w4001 = w4011 & w4050;
	assign w4000 = w4021 & w4040;
	assign w3944 = w4000 ^ w4001;
	assign w3999 = w4009 & w4041;
	assign w3994 = w4017 & w4049;
	assign w3993 = w4008 & w4053;
	assign w3960 = w4002 ^ w3993;
	assign w3992 = w4011 & w4046;
	assign w3962 = w4000 ^ w3992;
	assign w3991 = w4021 & w4047;
	assign w3990 = w4009 & w4052;
	assign w43701 = w4001 ^ w4002;
	assign w43703 = w4015 ^ w4033;
	assign w4007 = w43703 ^ w3985;
	assign w4005 = w4007 & w4044;
	assign w3996 = w4007 & w4048;
	assign w43702 = w4003 ^ w4005;
	assign w3974 = w25 ^ w43703;
	assign w4014 = w3974 ^ w3937;
	assign w3927 = w3974 ^ w3935;
	assign w3934 = w3964 ^ w3927;
	assign w4010 = w3931 ^ w3934;
	assign w4006 = w3927 ^ w3928;
	assign w4004 = w4014 & w4043;
	assign w3998 = w4006 & w4039;
	assign w3983 = w3998 ^ w43701;
	assign w3959 = w3998 ^ w4001;
	assign w3956 = ~w3959;
	assign w3955 = w3998 ^ w3999;
	assign w3949 = w3994 ^ w3983;
	assign w3946 = ~w3949;
	assign w3943 = w3999 ^ w3983;
	assign w3997 = w4010 & w4042;
	assign w3975 = w3993 ^ w3997;
	assign w3953 = ~w3975;
	assign w3952 = w3953 ^ w3991;
	assign w3948 = w3952 ^ w43702;
	assign w3951 = w3990 ^ w3948;
	assign w3995 = w4014 & w4045;
	assign w3989 = w4006 & w4054;
	assign w3988 = w4010 & w4051;
	assign w3954 = w3999 ^ w3988;
	assign w3950 = ~w3954;
	assign w4055 = w3950 ^ w3951;
	assign w47898 = ~w4055;
	assign w1888 = w229 ^ w47898;
	assign w1919 = w197 ^ w1888;
	assign w1951 = w165 ^ w1919;
	assign w1983 = w133 ^ w1951;
	assign w43517 = w3989 ^ w3990;
	assign w3958 = w3962 ^ w43517;
	assign w3961 = w43702 ^ w3958;
	assign w4058 = w3960 ^ w3961;
	assign w3957 = w3953 ^ w3958;
	assign w4057 = w3956 ^ w3957;
	assign w47893 = ~w4058;
	assign w1883 = w224 ^ w47893;
	assign w1914 = w192 ^ w1883;
	assign w1946 = w160 ^ w1914;
	assign w47894 = ~w4057;
	assign w1884 = w225 ^ w47894;
	assign w1915 = w193 ^ w1884;
	assign w1947 = w161 ^ w1915;
	assign w1979 = w129 ^ w1947;
	assign w1978 = w128 ^ w1946;
	assign w3971 = w3995 ^ w43517;
	assign w3972 = w3996 ^ w3971;
	assign w3976 = w4004 ^ w3972;
	assign w3981 = w4005 ^ w3976;
	assign w47897 = w43701 ^ w3981;
	assign w1887 = w228 ^ w47897;
	assign w1918 = w196 ^ w1887;
	assign w4056 = w3981 ^ w3955;
	assign w3947 = w3971 ^ w3948;
	assign w47895 = w3946 ^ w3947;
	assign w1885 = w226 ^ w47895;
	assign w1916 = w194 ^ w1885;
	assign w1948 = w162 ^ w1916;
	assign w3945 = w4003 ^ w3976;
	assign w47896 = w3944 ^ w3945;
	assign w1886 = w227 ^ w47896;
	assign w1917 = w195 ^ w1886;
	assign w1949 = w163 ^ w1917;
	assign w47900 = w3972 ^ w3943;
	assign w1890 = w231 ^ w47900;
	assign w1921 = w199 ^ w1890;
	assign w1953 = w167 ^ w1921;
	assign w1950 = w164 ^ w1918;
	assign w47899 = ~w4056;
	assign w1889 = w230 ^ w47899;
	assign w1920 = w198 ^ w1889;
	assign w1952 = w166 ^ w1920;
	assign w1984 = w134 ^ w1952;
	assign w4507 = w1978 ^ w1984;
	assign w4587 = w1983 ^ w4507;
	assign w4583 = w1979 ^ w4587;
	assign w4570 = w4587 & w4583;
	assign w1985 = w135 ^ w1953;
	assign w4501 = w1983 ^ w1985;
	assign w4584 = w4501 ^ w4507;
	assign w4590 = w1985 ^ w1979;
	assign w1982 = w132 ^ w1950;
	assign w4503 = w1982 ^ w1984;
	assign w4589 = w1982 ^ w1985;
	assign w4463 = w4503 ^ w4501;
	assign w4462 = w4503 ^ w1983;
	assign w4586 = w1978 ^ w4462;
	assign w4572 = w4586 & w1978;
	assign w1981 = w131 ^ w1949;
	assign w4500 = w1979 ^ w1981;
	assign w4581 = w4500 ^ w4589;
	assign w4580 = w1978 ^ w4581;
	assign w4579 = w4500 ^ w4463;
	assign w1980 = w130 ^ w1948;
	assign w4502 = w1980 ^ w4500;
	assign w4578 = w1984 ^ w4502;
	assign w4575 = w1983 ^ w4502;
	assign w4577 = w4507 ^ w4502;
	assign w4517 = w1979 ^ w1980;
	assign w4582 = w4517 ^ w4584;
	assign w4585 = w4589 ^ w4517;
	assign w4591 = w1980 ^ w1982;
	assign w4576 = w4501 ^ w4591;
	assign w4477 = w1981 ^ w1980;
	assign w4588 = w1985 ^ w1980;
	assign w4574 = w4581 & w4585;
	assign w4506 = w4574 ^ w4503;
	assign w4573 = w4582 & w4580;
	assign w4571 = w4590 & w4575;
	assign w4505 = w4571 ^ w4501;
	assign w4569 = w4584 & w4577;
	assign w4568 = w4589 & w4578;
	assign w4504 = w4568 ^ w4502;
	assign w4510 = w4506 ^ w4504;
	assign w4515 = w1985 ^ w4510;
	assign w4567 = w4591 & w4576;
	assign w4524 = w4567 ^ w4573;
	assign w4565 = w4524 ^ w4515;
	assign w4476 = w4567 ^ w4568;
	assign w4523 = w4476 ^ w4477;
	assign w4522 = w4523 ^ w4505;
	assign w4564 = w4570 ^ w4522;
	assign w4566 = w4588 & w4579;
	assign w4561 = w4565 & w4564;
	assign w43709 = w4298 ^ w4301;
	assign w4211 = w4237 ^ w43709;
	assign w4295 = w4211 ^ w4236;
	assign w4292 = w4293 ^ w4295;
	assign w4251 = w4299 ^ w43709;
	assign w4207 = w4302 ^ w4251;
	assign w4289 = w1995 ^ w4207;
	assign w43712 = w4298 ^ w4304;
	assign w4210 = w4242 ^ w43712;
	assign w4253 = w1999 ^ w4210;
	assign w4288 = w4293 ^ w4253;
	assign w4287 = w4288 & w4289;
	assign w4286 = w4287 ^ w4295;
	assign w4285 = w4293 ^ w4287;
	assign w4206 = w4287 ^ w4251;
	assign w4205 = w4287 ^ w4304;
	assign w4200 = w4205 ^ w4301;
	assign w4284 = w4295 & w4285;
	assign w4282 = w4284 ^ w4292;
	assign w4272 = w4286 & w1994;
	assign w4263 = w4286 & w4318;
	assign w43711 = w4284 ^ w4302;
	assign w4276 = w43711 ^ w4254;
	assign w4274 = w4276 & w4313;
	assign w4265 = w4276 & w4317;
	assign w4243 = w1995 ^ w43711;
	assign w4283 = w4243 ^ w4206;
	assign w4273 = w4283 & w4312;
	assign w4264 = w4283 & w4314;
	assign w4248 = w43712 ^ w4233;
	assign w4294 = w4256 ^ w4248;
	assign w4291 = w4294 & w4292;
	assign w4290 = w4291 ^ w4253;
	assign w4202 = w4291 ^ w4303;
	assign w4198 = w4202 ^ w4238;
	assign w4201 = w2001 ^ w4198;
	assign w4278 = w4200 ^ w4201;
	assign w4199 = w4291 ^ w4247;
	assign w4197 = w1999 ^ w4198;
	assign w4281 = w4290 & w4282;
	assign w4246 = w4281 ^ w4256;
	assign w4280 = w4246 ^ w4248;
	assign w4204 = w4281 ^ w4305;
	assign w4196 = w4243 ^ w4204;
	assign w4203 = w4233 ^ w4196;
	assign w4279 = w4200 ^ w4203;
	assign w4277 = w4246 ^ w4199;
	assign w4275 = w4196 ^ w4197;
	assign w4271 = w4277 & w4307;
	assign w4270 = w4280 & w4319;
	assign w4269 = w4290 & w4309;
	assign w4213 = w4269 ^ w4270;
	assign w4268 = w4278 & w4310;
	assign w4267 = w4275 & w4308;
	assign w4228 = w4267 ^ w4270;
	assign w4225 = ~w4228;
	assign w4224 = w4267 ^ w4268;
	assign w4266 = w4279 & w4311;
	assign w4262 = w4277 & w4322;
	assign w4244 = w4262 ^ w4266;
	assign w4229 = w4271 ^ w4262;
	assign w4222 = ~w4244;
	assign w4261 = w4280 & w4315;
	assign w4231 = w4269 ^ w4261;
	assign w4260 = w4290 & w4316;
	assign w4221 = w4222 ^ w4260;
	assign w4259 = w4278 & w4321;
	assign w4258 = w4275 & w4323;
	assign w4257 = w4279 & w4320;
	assign w4223 = w4268 ^ w4257;
	assign w4219 = ~w4223;
	assign w43710 = w4258 ^ w4259;
	assign w4240 = w4264 ^ w43710;
	assign w4241 = w4265 ^ w4240;
	assign w4245 = w4273 ^ w4241;
	assign w4250 = w4274 ^ w4245;
	assign w4325 = w4250 ^ w4224;
	assign w4214 = w4272 ^ w4245;
	assign w47944 = w4213 ^ w4214;
	assign w47947 = ~w4325;
	assign w2029 = w115 ^ w47944;
	assign w2032 = w118 ^ w47947;
	assign w1395 = w86 ^ w2032;
	assign w1427 = w54 ^ w1395;
	assign w1392 = w83 ^ w2029;
	assign w1424 = w51 ^ w1392;
	assign w1459 = w22 ^ w1427;
	assign w1456 = w19 ^ w1424;
	assign w4227 = w4231 ^ w43710;
	assign w4226 = w4222 ^ w4227;
	assign w4326 = w4225 ^ w4226;
	assign w47942 = ~w4326;
	assign w2027 = w113 ^ w47942;
	assign w1390 = w81 ^ w2027;
	assign w1422 = w49 ^ w1390;
	assign w1454 = w17 ^ w1422;
	assign w4634 = w1454 ^ w1456;
	assign w43713 = w4270 ^ w4271;
	assign w47945 = w43713 ^ w4250;
	assign w2030 = w116 ^ w47945;
	assign w1393 = w84 ^ w2030;
	assign w1425 = w52 ^ w1393;
	assign w1457 = w20 ^ w1425;
	assign w4637 = w1457 ^ w1459;
	assign w4252 = w4267 ^ w43713;
	assign w4218 = w4263 ^ w4252;
	assign w4215 = ~w4218;
	assign w4212 = w4268 ^ w4252;
	assign w47948 = w4241 ^ w4212;
	assign w2033 = w119 ^ w47948;
	assign w1396 = w87 ^ w2033;
	assign w1428 = w55 ^ w1396;
	assign w1460 = w23 ^ w1428;
	assign w4723 = w1457 ^ w1460;
	assign w4715 = w4634 ^ w4723;
	assign w4724 = w1460 ^ w1454;
	assign w43714 = w4272 ^ w4274;
	assign w4230 = w43714 ^ w4227;
	assign w4327 = w4229 ^ w4230;
	assign w47941 = ~w4327;
	assign w2026 = w112 ^ w47941;
	assign w1389 = w80 ^ w2026;
	assign w1421 = w48 ^ w1389;
	assign w1453 = w16 ^ w1421;
	assign w4641 = w1453 ^ w1459;
	assign w4714 = w1453 ^ w4715;
	assign w4217 = w4221 ^ w43714;
	assign w4220 = w4259 ^ w4217;
	assign w4324 = w4219 ^ w4220;
	assign w4216 = w4240 ^ w4217;
	assign w47943 = w4215 ^ w4216;
	assign w47946 = ~w4324;
	assign w2031 = w117 ^ w47946;
	assign w2028 = w114 ^ w47943;
	assign w1391 = w82 ^ w2028;
	assign w1394 = w85 ^ w2031;
	assign w1426 = w53 ^ w1394;
	assign w1423 = w50 ^ w1391;
	assign w1458 = w21 ^ w1426;
	assign w4635 = w1458 ^ w1460;
	assign w4718 = w4635 ^ w4641;
	assign w4721 = w1458 ^ w4641;
	assign w4717 = w1454 ^ w4721;
	assign w4597 = w4637 ^ w4635;
	assign w4713 = w4634 ^ w4597;
	assign w4596 = w4637 ^ w1458;
	assign w4720 = w1453 ^ w4596;
	assign w4706 = w4720 & w1453;
	assign w4704 = w4721 & w4717;
	assign w1455 = w18 ^ w1423;
	assign w4636 = w1455 ^ w4634;
	assign w4712 = w1459 ^ w4636;
	assign w4709 = w1458 ^ w4636;
	assign w4711 = w4641 ^ w4636;
	assign w4651 = w1454 ^ w1455;
	assign w4716 = w4651 ^ w4718;
	assign w4719 = w4723 ^ w4651;
	assign w4725 = w1455 ^ w1457;
	assign w4710 = w4635 ^ w4725;
	assign w4611 = w1456 ^ w1455;
	assign w4722 = w1460 ^ w1455;
	assign w4708 = w4715 & w4719;
	assign w4640 = w4708 ^ w4637;
	assign w4707 = w4716 & w4714;
	assign w4705 = w4724 & w4709;
	assign w4639 = w4705 ^ w4635;
	assign w4703 = w4718 & w4711;
	assign w4702 = w4723 & w4712;
	assign w4638 = w4702 ^ w4636;
	assign w4644 = w4640 ^ w4638;
	assign w4649 = w1460 ^ w4644;
	assign w4701 = w4725 & w4710;
	assign w4658 = w4701 ^ w4707;
	assign w4699 = w4658 ^ w4649;
	assign w4610 = w4701 ^ w4702;
	assign w4657 = w4610 ^ w4611;
	assign w4656 = w4657 ^ w4639;
	assign w4698 = w4704 ^ w4656;
	assign w4700 = w4722 & w4713;
	assign w4695 = w4699 & w4698;
	assign w43715 = w4432 ^ w4438;
	assign w4382 = w43715 ^ w4367;
	assign w4428 = w4390 ^ w4382;
	assign w4344 = w4376 ^ w43715;
	assign w4387 = w1991 ^ w4344;
	assign w4422 = w4427 ^ w4387;
	assign w43716 = w4432 ^ w4435;
	assign w4385 = w4433 ^ w43716;
	assign w4341 = w4436 ^ w4385;
	assign w4423 = w1987 ^ w4341;
	assign w4421 = w4422 & w4423;
	assign w4419 = w4427 ^ w4421;
	assign w4340 = w4421 ^ w4385;
	assign w4339 = w4421 ^ w4438;
	assign w4334 = w4339 ^ w4435;
	assign w4345 = w4371 ^ w43716;
	assign w4429 = w4345 ^ w4370;
	assign w4420 = w4421 ^ w4429;
	assign w4426 = w4427 ^ w4429;
	assign w4425 = w4428 & w4426;
	assign w4424 = w4425 ^ w4387;
	assign w4336 = w4425 ^ w4437;
	assign w4332 = w4336 ^ w4372;
	assign w4335 = w1993 ^ w4332;
	assign w4412 = w4334 ^ w4335;
	assign w4333 = w4425 ^ w4381;
	assign w4331 = w1991 ^ w4332;
	assign w4418 = w4429 & w4419;
	assign w4416 = w4418 ^ w4426;
	assign w4415 = w4424 & w4416;
	assign w4380 = w4415 ^ w4390;
	assign w4414 = w4380 ^ w4382;
	assign w4338 = w4415 ^ w4439;
	assign w4411 = w4380 ^ w4333;
	assign w4406 = w4420 & w1986;
	assign w4405 = w4411 & w4441;
	assign w4404 = w4414 & w4453;
	assign w4403 = w4424 & w4443;
	assign w4347 = w4403 ^ w4404;
	assign w4402 = w4412 & w4444;
	assign w4397 = w4420 & w4452;
	assign w4396 = w4411 & w4456;
	assign w4363 = w4405 ^ w4396;
	assign w4395 = w4414 & w4449;
	assign w4365 = w4403 ^ w4395;
	assign w4394 = w4424 & w4450;
	assign w4393 = w4412 & w4455;
	assign w43717 = w4404 ^ w4405;
	assign w43719 = w4418 ^ w4436;
	assign w4377 = w1987 ^ w43719;
	assign w4417 = w4377 ^ w4340;
	assign w4330 = w4377 ^ w4338;
	assign w4337 = w4367 ^ w4330;
	assign w4413 = w4334 ^ w4337;
	assign w4409 = w4330 ^ w4331;
	assign w4407 = w4417 & w4446;
	assign w4401 = w4409 & w4442;
	assign w4362 = w4401 ^ w4404;
	assign w4359 = ~w4362;
	assign w4358 = w4401 ^ w4402;
	assign w4400 = w4413 & w4445;
	assign w4398 = w4417 & w4448;
	assign w4378 = w4396 ^ w4400;
	assign w4356 = ~w4378;
	assign w4355 = w4356 ^ w4394;
	assign w4392 = w4409 & w4457;
	assign w4391 = w4413 & w4454;
	assign w4357 = w4402 ^ w4391;
	assign w4353 = ~w4357;
	assign w43518 = w4392 ^ w4393;
	assign w4361 = w4365 ^ w43518;
	assign w4360 = w4356 ^ w4361;
	assign w4460 = w4359 ^ w4360;
	assign w47934 = ~w4460;
	assign w2019 = w105 ^ w47934;
	assign w1382 = w73 ^ w2019;
	assign w1414 = w41 ^ w1382;
	assign w1446 = w9 ^ w1414;
	assign w4374 = w4398 ^ w43518;
	assign w4386 = w4401 ^ w43717;
	assign w4352 = w4397 ^ w4386;
	assign w4349 = ~w4352;
	assign w4346 = w4402 ^ w4386;
	assign w4410 = w43719 ^ w4388;
	assign w4408 = w4410 & w4447;
	assign w4399 = w4410 & w4451;
	assign w4375 = w4399 ^ w4374;
	assign w4379 = w4407 ^ w4375;
	assign w4384 = w4408 ^ w4379;
	assign w47937 = w43717 ^ w4384;
	assign w4459 = w4384 ^ w4358;
	assign w4348 = w4406 ^ w4379;
	assign w47936 = w4347 ^ w4348;
	assign w47940 = w4375 ^ w4346;
	assign w47939 = ~w4459;
	assign w2025 = w111 ^ w47940;
	assign w2024 = w110 ^ w47939;
	assign w2021 = w107 ^ w47936;
	assign w2022 = w108 ^ w47937;
	assign w1388 = w79 ^ w2025;
	assign w1420 = w47 ^ w1388;
	assign w1387 = w78 ^ w2024;
	assign w1419 = w46 ^ w1387;
	assign w1385 = w76 ^ w2022;
	assign w1417 = w44 ^ w1385;
	assign w1384 = w75 ^ w2021;
	assign w1416 = w43 ^ w1384;
	assign w1448 = w11 ^ w1416;
	assign w1452 = w15 ^ w1420;
	assign w1451 = w14 ^ w1419;
	assign w1449 = w12 ^ w1417;
	assign w35761 = w1446 ^ w1448;
	assign w35764 = w1449 ^ w1451;
	assign w35850 = w1449 ^ w1452;
	assign w35842 = w35761 ^ w35850;
	assign w35851 = w1452 ^ w1446;
	assign w43718 = w4406 ^ w4408;
	assign w4364 = w43718 ^ w4361;
	assign w4461 = w4363 ^ w4364;
	assign w47933 = ~w4461;
	assign w2018 = w104 ^ w47933;
	assign w1381 = w72 ^ w2018;
	assign w1413 = w40 ^ w1381;
	assign w1445 = w8 ^ w1413;
	assign w35768 = w1445 ^ w1451;
	assign w35841 = w1445 ^ w35842;
	assign w4351 = w4355 ^ w43718;
	assign w4354 = w4393 ^ w4351;
	assign w4458 = w4353 ^ w4354;
	assign w4350 = w4374 ^ w4351;
	assign w47935 = w4349 ^ w4350;
	assign w47938 = ~w4458;
	assign w2020 = w106 ^ w47935;
	assign w2023 = w109 ^ w47938;
	assign w1386 = w77 ^ w2023;
	assign w1418 = w45 ^ w1386;
	assign w1383 = w74 ^ w2020;
	assign w1415 = w42 ^ w1383;
	assign w1450 = w13 ^ w1418;
	assign w1447 = w10 ^ w1415;
	assign w35762 = w1450 ^ w1452;
	assign w35763 = w1447 ^ w35761;
	assign w35839 = w1451 ^ w35763;
	assign w35836 = w1450 ^ w35763;
	assign w35838 = w35768 ^ w35763;
	assign w35845 = w35762 ^ w35768;
	assign w35778 = w1446 ^ w1447;
	assign w35843 = w35778 ^ w35845;
	assign w35846 = w35850 ^ w35778;
	assign w35852 = w1447 ^ w1449;
	assign w35837 = w35762 ^ w35852;
	assign w35848 = w1450 ^ w35768;
	assign w35844 = w1446 ^ w35848;
	assign w35738 = w1448 ^ w1447;
	assign w35724 = w35764 ^ w35762;
	assign w35840 = w35761 ^ w35724;
	assign w35723 = w35764 ^ w1450;
	assign w35847 = w1445 ^ w35723;
	assign w35849 = w1452 ^ w1447;
	assign w35835 = w35842 & w35846;
	assign w35767 = w35835 ^ w35764;
	assign w35834 = w35843 & w35841;
	assign w35833 = w35847 & w1445;
	assign w35832 = w35851 & w35836;
	assign w35766 = w35832 ^ w35762;
	assign w35831 = w35848 & w35844;
	assign w35830 = w35845 & w35838;
	assign w35829 = w35850 & w35839;
	assign w35765 = w35829 ^ w35763;
	assign w35771 = w35767 ^ w35765;
	assign w35776 = w1452 ^ w35771;
	assign w35828 = w35852 & w35837;
	assign w35785 = w35828 ^ w35834;
	assign w35826 = w35785 ^ w35776;
	assign w35737 = w35828 ^ w35829;
	assign w35784 = w35737 ^ w35738;
	assign w35783 = w35784 ^ w35766;
	assign w35825 = w35831 ^ w35783;
	assign w35827 = w35849 & w35840;
	assign w35822 = w35826 & w35825;
	assign w43720 = w4566 ^ w4572;
	assign w4478 = w4510 ^ w43720;
	assign w4521 = w1983 ^ w4478;
	assign w4556 = w4561 ^ w4521;
	assign w4516 = w43720 ^ w4501;
	assign w4562 = w4524 ^ w4516;
	assign w43721 = w4566 ^ w4569;
	assign w4519 = w4567 ^ w43721;
	assign w4475 = w4570 ^ w4519;
	assign w4557 = w1979 ^ w4475;
	assign w4555 = w4556 & w4557;
	assign w4553 = w4561 ^ w4555;
	assign w4474 = w4555 ^ w4519;
	assign w4473 = w4555 ^ w4572;
	assign w4468 = w4473 ^ w4569;
	assign w4479 = w4505 ^ w43721;
	assign w4563 = w4479 ^ w4504;
	assign w4554 = w4555 ^ w4563;
	assign w4560 = w4561 ^ w4563;
	assign w4559 = w4562 & w4560;
	assign w4558 = w4559 ^ w4521;
	assign w4470 = w4559 ^ w4571;
	assign w4466 = w4470 ^ w4506;
	assign w4469 = w1985 ^ w4466;
	assign w4546 = w4468 ^ w4469;
	assign w4467 = w4559 ^ w4515;
	assign w4465 = w1983 ^ w4466;
	assign w4552 = w4563 & w4553;
	assign w4550 = w4552 ^ w4560;
	assign w4549 = w4558 & w4550;
	assign w4514 = w4549 ^ w4524;
	assign w4548 = w4514 ^ w4516;
	assign w4472 = w4549 ^ w4573;
	assign w4545 = w4514 ^ w4467;
	assign w4540 = w4554 & w1978;
	assign w4539 = w4545 & w4575;
	assign w4538 = w4548 & w4587;
	assign w4537 = w4558 & w4577;
	assign w4481 = w4537 ^ w4538;
	assign w4536 = w4546 & w4578;
	assign w4531 = w4554 & w4586;
	assign w4530 = w4545 & w4590;
	assign w4497 = w4539 ^ w4530;
	assign w4529 = w4548 & w4583;
	assign w4499 = w4537 ^ w4529;
	assign w4528 = w4558 & w4584;
	assign w4527 = w4546 & w4589;
	assign w43723 = w4538 ^ w4539;
	assign w43725 = w4552 ^ w4570;
	assign w4544 = w43725 ^ w4522;
	assign w4542 = w4544 & w4581;
	assign w4533 = w4544 & w4585;
	assign w43724 = w4540 ^ w4542;
	assign w4511 = w1979 ^ w43725;
	assign w4551 = w4511 ^ w4474;
	assign w4464 = w4511 ^ w4472;
	assign w4471 = w4501 ^ w4464;
	assign w4547 = w4468 ^ w4471;
	assign w4543 = w4464 ^ w4465;
	assign w4541 = w4551 & w4580;
	assign w4535 = w4543 & w4576;
	assign w4520 = w4535 ^ w43723;
	assign w4496 = w4535 ^ w4538;
	assign w4493 = ~w4496;
	assign w4492 = w4535 ^ w4536;
	assign w4486 = w4531 ^ w4520;
	assign w4483 = ~w4486;
	assign w4480 = w4536 ^ w4520;
	assign w4534 = w4547 & w4579;
	assign w4512 = w4530 ^ w4534;
	assign w4490 = ~w4512;
	assign w4489 = w4490 ^ w4528;
	assign w4485 = w4489 ^ w43724;
	assign w4488 = w4527 ^ w4485;
	assign w4532 = w4551 & w4582;
	assign w4526 = w4543 & w4591;
	assign w4525 = w4547 & w4588;
	assign w4491 = w4536 ^ w4525;
	assign w4487 = ~w4491;
	assign w4592 = w4487 ^ w4488;
	assign w47930 = ~w4592;
	assign w2015 = w101 ^ w47930;
	assign w1378 = w69 ^ w2015;
	assign w1410 = w37 ^ w1378;
	assign w1442 = w5 ^ w1410;
	assign w43722 = w4526 ^ w4527;
	assign w4495 = w4499 ^ w43722;
	assign w4498 = w43724 ^ w4495;
	assign w4595 = w4497 ^ w4498;
	assign w4494 = w4490 ^ w4495;
	assign w4594 = w4493 ^ w4494;
	assign w47925 = ~w4595;
	assign w47926 = ~w4594;
	assign w2011 = w97 ^ w47926;
	assign w2010 = w96 ^ w47925;
	assign w1373 = w64 ^ w2010;
	assign w1374 = w65 ^ w2011;
	assign w1406 = w33 ^ w1374;
	assign w1405 = w32 ^ w1373;
	assign w1438 = w1 ^ w1406;
	assign w1437 = w0 ^ w1405;
	assign w4508 = w4532 ^ w43722;
	assign w4509 = w4533 ^ w4508;
	assign w4513 = w4541 ^ w4509;
	assign w4518 = w4542 ^ w4513;
	assign w47929 = w43723 ^ w4518;
	assign w4593 = w4518 ^ w4492;
	assign w4484 = w4508 ^ w4485;
	assign w47927 = w4483 ^ w4484;
	assign w4482 = w4540 ^ w4513;
	assign w47928 = w4481 ^ w4482;
	assign w47932 = w4509 ^ w4480;
	assign w47931 = ~w4593;
	assign w2017 = w103 ^ w47932;
	assign w2016 = w102 ^ w47931;
	assign w2014 = w100 ^ w47929;
	assign w2013 = w99 ^ w47928;
	assign w2012 = w98 ^ w47927;
	assign w1377 = w68 ^ w2014;
	assign w1380 = w71 ^ w2017;
	assign w1412 = w39 ^ w1380;
	assign w1379 = w70 ^ w2016;
	assign w1376 = w67 ^ w2013;
	assign w1375 = w66 ^ w2012;
	assign w1408 = w35 ^ w1376;
	assign w1407 = w34 ^ w1375;
	assign w1411 = w38 ^ w1379;
	assign w1409 = w36 ^ w1377;
	assign w1440 = w3 ^ w1408;
	assign w1444 = w7 ^ w1412;
	assign w1439 = w2 ^ w1407;
	assign w1443 = w6 ^ w1411;
	assign w1441 = w4 ^ w1409;
	assign w23299 = w1438 ^ w1440;
	assign w23300 = w1442 ^ w1444;
	assign w23301 = w1439 ^ w23299;
	assign w23377 = w1443 ^ w23301;
	assign w23374 = w1442 ^ w23301;
	assign w23302 = w1441 ^ w1443;
	assign w23306 = w1437 ^ w1443;
	assign w23376 = w23306 ^ w23301;
	assign w23388 = w1441 ^ w1444;
	assign w23383 = w23300 ^ w23306;
	assign w23380 = w23299 ^ w23388;
	assign w23379 = w1437 ^ w23380;
	assign w23316 = w1438 ^ w1439;
	assign w23381 = w23316 ^ w23383;
	assign w23384 = w23388 ^ w23316;
	assign w23390 = w1439 ^ w1441;
	assign w23375 = w23300 ^ w23390;
	assign w23386 = w1442 ^ w23306;
	assign w23382 = w1438 ^ w23386;
	assign w23276 = w1440 ^ w1439;
	assign w23262 = w23302 ^ w23300;
	assign w23378 = w23299 ^ w23262;
	assign w23261 = w23302 ^ w1442;
	assign w23385 = w1437 ^ w23261;
	assign w23389 = w1444 ^ w1438;
	assign w23387 = w1444 ^ w1439;
	assign w23373 = w23380 & w23384;
	assign w23305 = w23373 ^ w23302;
	assign w23372 = w23381 & w23379;
	assign w23371 = w23385 & w1437;
	assign w23370 = w23389 & w23374;
	assign w23304 = w23370 ^ w23300;
	assign w23369 = w23386 & w23382;
	assign w23368 = w23383 & w23376;
	assign w23367 = w23388 & w23377;
	assign w23303 = w23367 ^ w23301;
	assign w23309 = w23305 ^ w23303;
	assign w23314 = w1444 ^ w23309;
	assign w23366 = w23390 & w23375;
	assign w23323 = w23366 ^ w23372;
	assign w23364 = w23323 ^ w23314;
	assign w23275 = w23366 ^ w23367;
	assign w23322 = w23275 ^ w23276;
	assign w23321 = w23322 ^ w23304;
	assign w23363 = w23369 ^ w23321;
	assign w23365 = w23387 & w23378;
	assign w23360 = w23364 & w23363;
	assign w43726 = w4700 ^ w4703;
	assign w4613 = w4639 ^ w43726;
	assign w4697 = w4613 ^ w4638;
	assign w4694 = w4695 ^ w4697;
	assign w4653 = w4701 ^ w43726;
	assign w4609 = w4704 ^ w4653;
	assign w4691 = w1454 ^ w4609;
	assign w43729 = w4700 ^ w4706;
	assign w4612 = w4644 ^ w43729;
	assign w4655 = w1458 ^ w4612;
	assign w4690 = w4695 ^ w4655;
	assign w4689 = w4690 & w4691;
	assign w4688 = w4689 ^ w4697;
	assign w4687 = w4695 ^ w4689;
	assign w4608 = w4689 ^ w4653;
	assign w4607 = w4689 ^ w4706;
	assign w4602 = w4607 ^ w4703;
	assign w4686 = w4697 & w4687;
	assign w4684 = w4686 ^ w4694;
	assign w4674 = w4688 & w1453;
	assign w4665 = w4688 & w4720;
	assign w43728 = w4686 ^ w4704;
	assign w4678 = w43728 ^ w4656;
	assign w4676 = w4678 & w4715;
	assign w4667 = w4678 & w4719;
	assign w4645 = w1454 ^ w43728;
	assign w4685 = w4645 ^ w4608;
	assign w4675 = w4685 & w4714;
	assign w4666 = w4685 & w4716;
	assign w4650 = w43729 ^ w4635;
	assign w4696 = w4658 ^ w4650;
	assign w4693 = w4696 & w4694;
	assign w4692 = w4693 ^ w4655;
	assign w4604 = w4693 ^ w4705;
	assign w4600 = w4604 ^ w4640;
	assign w4603 = w1460 ^ w4600;
	assign w4680 = w4602 ^ w4603;
	assign w4601 = w4693 ^ w4649;
	assign w4599 = w1458 ^ w4600;
	assign w4683 = w4692 & w4684;
	assign w4648 = w4683 ^ w4658;
	assign w4682 = w4648 ^ w4650;
	assign w4606 = w4683 ^ w4707;
	assign w4598 = w4645 ^ w4606;
	assign w4605 = w4635 ^ w4598;
	assign w4681 = w4602 ^ w4605;
	assign w4679 = w4648 ^ w4601;
	assign w4677 = w4598 ^ w4599;
	assign w4673 = w4679 & w4709;
	assign w4672 = w4682 & w4721;
	assign w4671 = w4692 & w4711;
	assign w4615 = w4671 ^ w4672;
	assign w4670 = w4680 & w4712;
	assign w4669 = w4677 & w4710;
	assign w4630 = w4669 ^ w4672;
	assign w4627 = ~w4630;
	assign w4626 = w4669 ^ w4670;
	assign w4668 = w4681 & w4713;
	assign w4664 = w4679 & w4724;
	assign w4646 = w4664 ^ w4668;
	assign w4631 = w4673 ^ w4664;
	assign w4624 = ~w4646;
	assign w4663 = w4682 & w4717;
	assign w4633 = w4671 ^ w4663;
	assign w4662 = w4692 & w4718;
	assign w4623 = w4624 ^ w4662;
	assign w4661 = w4680 & w4723;
	assign w4660 = w4677 & w4725;
	assign w4659 = w4681 & w4722;
	assign w4625 = w4670 ^ w4659;
	assign w4621 = ~w4625;
	assign w43727 = w4660 ^ w4661;
	assign w4642 = w4666 ^ w43727;
	assign w4643 = w4667 ^ w4642;
	assign w4647 = w4675 ^ w4643;
	assign w4652 = w4676 ^ w4647;
	assign w4727 = w4652 ^ w4626;
	assign w4616 = w4674 ^ w4647;
	assign w47984 = w4615 ^ w4616;
	assign w47987 = ~w4727;
	assign w1498 = w1912 ^ w47987;
	assign w1495 = w1909 ^ w47984;
	assign w1530 = w1944 ^ w1498;
	assign w1562 = w1976 ^ w1530;
	assign w1527 = w1941 ^ w1495;
	assign w1559 = w1973 ^ w1527;
	assign w1594 = w2008 ^ w1562;
	assign w1591 = w2005 ^ w1559;
	assign w4629 = w4633 ^ w43727;
	assign w4628 = w4624 ^ w4629;
	assign w4728 = w4627 ^ w4628;
	assign w47982 = ~w4728;
	assign w2043 = w1907 ^ w47982;
	assign w43730 = w4672 ^ w4673;
	assign w47985 = w43730 ^ w4652;
	assign w1496 = w1910 ^ w47985;
	assign w1528 = w1942 ^ w1496;
	assign w1560 = w1974 ^ w1528;
	assign w1592 = w2006 ^ w1560;
	assign w38444 = w1592 ^ w1594;
	assign w4654 = w4669 ^ w43730;
	assign w4620 = w4665 ^ w4654;
	assign w4617 = ~w4620;
	assign w4614 = w4670 ^ w4654;
	assign w47988 = w4643 ^ w4614;
	assign w1499 = w1913 ^ w47988;
	assign w1531 = w1945 ^ w1499;
	assign w1563 = w1977 ^ w1531;
	assign w1595 = w2009 ^ w1563;
	assign w38530 = w1592 ^ w1595;
	assign w43731 = w4674 ^ w4676;
	assign w4632 = w43731 ^ w4629;
	assign w4729 = w4631 ^ w4632;
	assign w47981 = ~w4729;
	assign w4619 = w4623 ^ w43731;
	assign w4622 = w4661 ^ w4619;
	assign w4726 = w4621 ^ w4622;
	assign w4618 = w4642 ^ w4619;
	assign w47983 = w4617 ^ w4618;
	assign w47986 = ~w4726;
	assign w1497 = w1911 ^ w47986;
	assign w1494 = w1908 ^ w47983;
	assign w1529 = w1943 ^ w1497;
	assign w1561 = w1975 ^ w1529;
	assign w1526 = w1940 ^ w1494;
	assign w1558 = w1972 ^ w1526;
	assign w1593 = w2007 ^ w1561;
	assign w1590 = w2004 ^ w1558;
	assign w38442 = w1593 ^ w1595;
	assign w38532 = w1590 ^ w1592;
	assign w38517 = w38442 ^ w38532;
	assign w38418 = w1591 ^ w1590;
	assign w38404 = w38444 ^ w38442;
	assign w38403 = w38444 ^ w1593;
	assign w38529 = w1595 ^ w1590;
	assign w38508 = w38532 & w38517;
	assign w43746 = w5238 ^ w5241;
	assign w5151 = w5177 ^ w43746;
	assign w5235 = w5151 ^ w5176;
	assign w5232 = w5233 ^ w5235;
	assign w5191 = w5239 ^ w43746;
	assign w5147 = w5242 ^ w5191;
	assign w5229 = w47883 ^ w5147;
	assign w43749 = w5238 ^ w5244;
	assign w5150 = w5182 ^ w43749;
	assign w5193 = w47879 ^ w5150;
	assign w5228 = w5233 ^ w5193;
	assign w5227 = w5228 & w5229;
	assign w5226 = w5227 ^ w5235;
	assign w5225 = w5233 ^ w5227;
	assign w5146 = w5227 ^ w5191;
	assign w5145 = w5227 ^ w5244;
	assign w5140 = w5145 ^ w5241;
	assign w5224 = w5235 & w5225;
	assign w5222 = w5224 ^ w5232;
	assign w5212 = w5226 & w47884;
	assign w5203 = w5226 & w5258;
	assign w43748 = w5224 ^ w5242;
	assign w5216 = w43748 ^ w5194;
	assign w5214 = w5216 & w5253;
	assign w5205 = w5216 & w5257;
	assign w5183 = w47883 ^ w43748;
	assign w5223 = w5183 ^ w5146;
	assign w5213 = w5223 & w5252;
	assign w5204 = w5223 & w5254;
	assign w5188 = w43749 ^ w5173;
	assign w5234 = w5196 ^ w5188;
	assign w5231 = w5234 & w5232;
	assign w5230 = w5231 ^ w5193;
	assign w5142 = w5231 ^ w5243;
	assign w5138 = w5142 ^ w5178;
	assign w5141 = w47877 ^ w5138;
	assign w5218 = w5140 ^ w5141;
	assign w5139 = w5231 ^ w5187;
	assign w5137 = w47879 ^ w5138;
	assign w5221 = w5230 & w5222;
	assign w5186 = w5221 ^ w5196;
	assign w5220 = w5186 ^ w5188;
	assign w5144 = w5221 ^ w5245;
	assign w5136 = w5183 ^ w5144;
	assign w5143 = w5173 ^ w5136;
	assign w5219 = w5140 ^ w5143;
	assign w5217 = w5186 ^ w5139;
	assign w5215 = w5136 ^ w5137;
	assign w5211 = w5217 & w5247;
	assign w5210 = w5220 & w5259;
	assign w5209 = w5230 & w5249;
	assign w5153 = w5209 ^ w5210;
	assign w5208 = w5218 & w5250;
	assign w5207 = w5215 & w5248;
	assign w5168 = w5207 ^ w5210;
	assign w5165 = ~w5168;
	assign w5164 = w5207 ^ w5208;
	assign w5206 = w5219 & w5251;
	assign w5202 = w5217 & w5262;
	assign w5184 = w5202 ^ w5206;
	assign w5169 = w5211 ^ w5202;
	assign w5162 = ~w5184;
	assign w5201 = w5220 & w5255;
	assign w5171 = w5209 ^ w5201;
	assign w5200 = w5230 & w5256;
	assign w5161 = w5162 ^ w5200;
	assign w5199 = w5218 & w5261;
	assign w5198 = w5215 & w5263;
	assign w5197 = w5219 & w5260;
	assign w5163 = w5208 ^ w5197;
	assign w5159 = ~w5163;
	assign w43747 = w5198 ^ w5199;
	assign w5180 = w5204 ^ w43747;
	assign w5181 = w5205 ^ w5180;
	assign w5185 = w5213 ^ w5181;
	assign w5190 = w5214 ^ w5185;
	assign w5265 = w5190 ^ w5164;
	assign w5154 = w5212 ^ w5185;
	assign w48480 = w5153 ^ w5154;
	assign w48483 = ~w5265;
	assign w6252 = ~w48480;
	assign w5167 = w5171 ^ w43747;
	assign w5166 = w5162 ^ w5167;
	assign w5266 = w5165 ^ w5166;
	assign w48478 = ~w5266;
	assign w43750 = w5210 ^ w5211;
	assign w48481 = w43750 ^ w5190;
	assign w5192 = w5207 ^ w43750;
	assign w5158 = w5203 ^ w5192;
	assign w5155 = ~w5158;
	assign w5152 = w5208 ^ w5192;
	assign w48484 = w5181 ^ w5152;
	assign w43751 = w5212 ^ w5214;
	assign w5170 = w43751 ^ w5167;
	assign w5267 = w5169 ^ w5170;
	assign w5157 = w5161 ^ w43751;
	assign w5160 = w5199 ^ w5157;
	assign w5264 = w5159 ^ w5160;
	assign w5156 = w5180 ^ w5157;
	assign w48479 = w5155 ^ w5156;
	assign w48482 = ~w5264;
	assign w6245 = ~w48479;
	assign w43752 = w5372 ^ w5375;
	assign w5285 = w5311 ^ w43752;
	assign w5369 = w5285 ^ w5310;
	assign w5366 = w5367 ^ w5369;
	assign w5325 = w5373 ^ w43752;
	assign w5281 = w5376 ^ w5325;
	assign w5363 = w47875 ^ w5281;
	assign w43755 = w5372 ^ w5378;
	assign w5284 = w5316 ^ w43755;
	assign w5327 = w47871 ^ w5284;
	assign w5362 = w5367 ^ w5327;
	assign w5361 = w5362 & w5363;
	assign w5360 = w5361 ^ w5369;
	assign w5359 = w5367 ^ w5361;
	assign w5280 = w5361 ^ w5325;
	assign w5279 = w5361 ^ w5378;
	assign w5274 = w5279 ^ w5375;
	assign w5358 = w5369 & w5359;
	assign w5356 = w5358 ^ w5366;
	assign w5346 = w5360 & w47876;
	assign w5337 = w5360 & w5392;
	assign w43754 = w5358 ^ w5376;
	assign w5350 = w43754 ^ w5328;
	assign w5348 = w5350 & w5387;
	assign w5339 = w5350 & w5391;
	assign w5317 = w47875 ^ w43754;
	assign w5357 = w5317 ^ w5280;
	assign w5347 = w5357 & w5386;
	assign w5338 = w5357 & w5388;
	assign w5322 = w43755 ^ w5307;
	assign w5368 = w5330 ^ w5322;
	assign w5365 = w5368 & w5366;
	assign w5364 = w5365 ^ w5327;
	assign w5276 = w5365 ^ w5377;
	assign w5272 = w5276 ^ w5312;
	assign w5275 = w47869 ^ w5272;
	assign w5352 = w5274 ^ w5275;
	assign w5273 = w5365 ^ w5321;
	assign w5271 = w47871 ^ w5272;
	assign w5355 = w5364 & w5356;
	assign w5320 = w5355 ^ w5330;
	assign w5354 = w5320 ^ w5322;
	assign w5278 = w5355 ^ w5379;
	assign w5270 = w5317 ^ w5278;
	assign w5277 = w5307 ^ w5270;
	assign w5353 = w5274 ^ w5277;
	assign w5351 = w5320 ^ w5273;
	assign w5349 = w5270 ^ w5271;
	assign w5345 = w5351 & w5381;
	assign w5344 = w5354 & w5393;
	assign w5343 = w5364 & w5383;
	assign w5287 = w5343 ^ w5344;
	assign w5342 = w5352 & w5384;
	assign w5341 = w5349 & w5382;
	assign w5302 = w5341 ^ w5344;
	assign w5299 = ~w5302;
	assign w5298 = w5341 ^ w5342;
	assign w5340 = w5353 & w5385;
	assign w5336 = w5351 & w5396;
	assign w5318 = w5336 ^ w5340;
	assign w5303 = w5345 ^ w5336;
	assign w5296 = ~w5318;
	assign w5335 = w5354 & w5389;
	assign w5305 = w5343 ^ w5335;
	assign w5334 = w5364 & w5390;
	assign w5295 = w5296 ^ w5334;
	assign w5333 = w5352 & w5395;
	assign w5332 = w5349 & w5397;
	assign w5331 = w5353 & w5394;
	assign w5297 = w5342 ^ w5331;
	assign w5293 = ~w5297;
	assign w43753 = w5332 ^ w5333;
	assign w5314 = w5338 ^ w43753;
	assign w5315 = w5339 ^ w5314;
	assign w5319 = w5347 ^ w5315;
	assign w5324 = w5348 ^ w5319;
	assign w5399 = w5324 ^ w5298;
	assign w5288 = w5346 ^ w5319;
	assign w48467 = w5287 ^ w5288;
	assign w5301 = w5305 ^ w43753;
	assign w5300 = w5296 ^ w5301;
	assign w5400 = w5299 ^ w5300;
	assign w43756 = w5344 ^ w5345;
	assign w48468 = w43756 ^ w5324;
	assign w6161 = ~w48468;
	assign w5326 = w5341 ^ w43756;
	assign w5292 = w5337 ^ w5326;
	assign w5289 = ~w5292;
	assign w5286 = w5342 ^ w5326;
	assign w48469 = w5315 ^ w5286;
	assign w43757 = w5346 ^ w5348;
	assign w5304 = w43757 ^ w5301;
	assign w5401 = w5303 ^ w5304;
	assign w5291 = w5295 ^ w43757;
	assign w5294 = w5333 ^ w5291;
	assign w5398 = w5293 ^ w5294;
	assign w5290 = w5314 ^ w5291;
	assign w48466 = w5289 ^ w5290;
	assign w43758 = w5506 ^ w5512;
	assign w5456 = w43758 ^ w5441;
	assign w5502 = w5464 ^ w5456;
	assign w5418 = w5450 ^ w43758;
	assign w5461 = w47863 ^ w5418;
	assign w5496 = w5501 ^ w5461;
	assign w43759 = w5506 ^ w5509;
	assign w5459 = w5507 ^ w43759;
	assign w5415 = w5510 ^ w5459;
	assign w5497 = w47867 ^ w5415;
	assign w5495 = w5496 & w5497;
	assign w5493 = w5501 ^ w5495;
	assign w5414 = w5495 ^ w5459;
	assign w5413 = w5495 ^ w5512;
	assign w5408 = w5413 ^ w5509;
	assign w5419 = w5445 ^ w43759;
	assign w5503 = w5419 ^ w5444;
	assign w5494 = w5495 ^ w5503;
	assign w5500 = w5501 ^ w5503;
	assign w5499 = w5502 & w5500;
	assign w5498 = w5499 ^ w5461;
	assign w5410 = w5499 ^ w5511;
	assign w5406 = w5410 ^ w5446;
	assign w5409 = w47861 ^ w5406;
	assign w5486 = w5408 ^ w5409;
	assign w5407 = w5499 ^ w5455;
	assign w5405 = w47863 ^ w5406;
	assign w5492 = w5503 & w5493;
	assign w5490 = w5492 ^ w5500;
	assign w5489 = w5498 & w5490;
	assign w5454 = w5489 ^ w5464;
	assign w5488 = w5454 ^ w5456;
	assign w5412 = w5489 ^ w5513;
	assign w5485 = w5454 ^ w5407;
	assign w5480 = w5494 & w47868;
	assign w5479 = w5485 & w5515;
	assign w5478 = w5488 & w5527;
	assign w5477 = w5498 & w5517;
	assign w5421 = w5477 ^ w5478;
	assign w5476 = w5486 & w5518;
	assign w5471 = w5494 & w5526;
	assign w5470 = w5485 & w5530;
	assign w5437 = w5479 ^ w5470;
	assign w5469 = w5488 & w5523;
	assign w5439 = w5477 ^ w5469;
	assign w5468 = w5498 & w5524;
	assign w5467 = w5486 & w5529;
	assign w43760 = w5478 ^ w5479;
	assign w43762 = w5492 ^ w5510;
	assign w5451 = w47867 ^ w43762;
	assign w5491 = w5451 ^ w5414;
	assign w5404 = w5451 ^ w5412;
	assign w5411 = w5441 ^ w5404;
	assign w5487 = w5408 ^ w5411;
	assign w5483 = w5404 ^ w5405;
	assign w5481 = w5491 & w5520;
	assign w5475 = w5483 & w5516;
	assign w5436 = w5475 ^ w5478;
	assign w5433 = ~w5436;
	assign w5432 = w5475 ^ w5476;
	assign w5474 = w5487 & w5519;
	assign w5472 = w5491 & w5522;
	assign w5452 = w5470 ^ w5474;
	assign w5430 = ~w5452;
	assign w5429 = w5430 ^ w5468;
	assign w5466 = w5483 & w5531;
	assign w5465 = w5487 & w5528;
	assign w5431 = w5476 ^ w5465;
	assign w5427 = ~w5431;
	assign w43521 = w5466 ^ w5467;
	assign w5448 = w5472 ^ w43521;
	assign w5435 = w5439 ^ w43521;
	assign w5434 = w5430 ^ w5435;
	assign w5534 = w5433 ^ w5434;
	assign w5460 = w5475 ^ w43760;
	assign w5426 = w5471 ^ w5460;
	assign w5423 = ~w5426;
	assign w5420 = w5476 ^ w5460;
	assign w5484 = w43762 ^ w5462;
	assign w5482 = w5484 & w5521;
	assign w5473 = w5484 & w5525;
	assign w5449 = w5473 ^ w5448;
	assign w5453 = w5481 ^ w5449;
	assign w5458 = w5482 ^ w5453;
	assign w48454 = w43760 ^ w5458;
	assign w5533 = w5458 ^ w5432;
	assign w5422 = w5480 ^ w5453;
	assign w48453 = w5421 ^ w5422;
	assign w48456 = w5449 ^ w5420;
	assign w48455 = ~w5533;
	assign w43761 = w5480 ^ w5482;
	assign w5438 = w43761 ^ w5435;
	assign w5535 = w5437 ^ w5438;
	assign w5425 = w5429 ^ w43761;
	assign w5428 = w5467 ^ w5425;
	assign w5532 = w5427 ^ w5428;
	assign w5424 = w5448 ^ w5425;
	assign w48452 = w5423 ^ w5424;
	assign w43763 = w5640 ^ w5646;
	assign w5552 = w5584 ^ w43763;
	assign w5595 = w47847 ^ w5552;
	assign w5630 = w5635 ^ w5595;
	assign w5590 = w43763 ^ w5575;
	assign w5636 = w5598 ^ w5590;
	assign w43764 = w5640 ^ w5643;
	assign w5593 = w5641 ^ w43764;
	assign w5549 = w5644 ^ w5593;
	assign w5631 = w47851 ^ w5549;
	assign w5629 = w5630 & w5631;
	assign w5548 = w5629 ^ w5593;
	assign w5547 = w5629 ^ w5646;
	assign w5542 = w5547 ^ w5643;
	assign w5627 = w5635 ^ w5629;
	assign w5553 = w5579 ^ w43764;
	assign w5637 = w5553 ^ w5578;
	assign w5628 = w5629 ^ w5637;
	assign w5634 = w5635 ^ w5637;
	assign w5633 = w5636 & w5634;
	assign w5632 = w5633 ^ w5595;
	assign w5544 = w5633 ^ w5645;
	assign w5540 = w5544 ^ w5580;
	assign w5543 = w47845 ^ w5540;
	assign w5620 = w5542 ^ w5543;
	assign w5541 = w5633 ^ w5589;
	assign w5539 = w47847 ^ w5540;
	assign w5626 = w5637 & w5627;
	assign w5624 = w5626 ^ w5634;
	assign w5623 = w5632 & w5624;
	assign w5588 = w5623 ^ w5598;
	assign w5622 = w5588 ^ w5590;
	assign w5546 = w5623 ^ w5647;
	assign w5619 = w5588 ^ w5541;
	assign w5614 = w5628 & w47852;
	assign w5613 = w5619 & w5649;
	assign w5612 = w5622 & w5661;
	assign w5611 = w5632 & w5651;
	assign w5555 = w5611 ^ w5612;
	assign w5610 = w5620 & w5652;
	assign w5605 = w5628 & w5660;
	assign w5604 = w5619 & w5664;
	assign w5571 = w5613 ^ w5604;
	assign w5603 = w5622 & w5657;
	assign w5573 = w5611 ^ w5603;
	assign w5602 = w5632 & w5658;
	assign w5601 = w5620 & w5663;
	assign w43766 = w5612 ^ w5613;
	assign w43768 = w5626 ^ w5644;
	assign w5618 = w43768 ^ w5596;
	assign w5616 = w5618 & w5655;
	assign w5607 = w5618 & w5659;
	assign w43767 = w5614 ^ w5616;
	assign w5585 = w47851 ^ w43768;
	assign w5625 = w5585 ^ w5548;
	assign w5538 = w5585 ^ w5546;
	assign w5545 = w5575 ^ w5538;
	assign w5621 = w5542 ^ w5545;
	assign w5617 = w5538 ^ w5539;
	assign w5615 = w5625 & w5654;
	assign w5609 = w5617 & w5650;
	assign w5594 = w5609 ^ w43766;
	assign w5570 = w5609 ^ w5612;
	assign w5567 = ~w5570;
	assign w5566 = w5609 ^ w5610;
	assign w5560 = w5605 ^ w5594;
	assign w5557 = ~w5560;
	assign w5554 = w5610 ^ w5594;
	assign w5608 = w5621 & w5653;
	assign w5586 = w5604 ^ w5608;
	assign w5564 = ~w5586;
	assign w5563 = w5564 ^ w5602;
	assign w5559 = w5563 ^ w43767;
	assign w5562 = w5601 ^ w5559;
	assign w5606 = w5625 & w5656;
	assign w5600 = w5617 & w5665;
	assign w5599 = w5621 & w5662;
	assign w5565 = w5610 ^ w5599;
	assign w5561 = ~w5565;
	assign w5666 = w5561 ^ w5562;
	assign w43765 = w5600 ^ w5601;
	assign w5582 = w5606 ^ w43765;
	assign w5583 = w5607 ^ w5582;
	assign w5587 = w5615 ^ w5583;
	assign w5592 = w5616 ^ w5587;
	assign w48500 = w43766 ^ w5592;
	assign w5667 = w5592 ^ w5566;
	assign w5558 = w5582 ^ w5559;
	assign w48498 = w5557 ^ w5558;
	assign w5556 = w5614 ^ w5587;
	assign w48499 = w5555 ^ w5556;
	assign w48501 = w5583 ^ w5554;
	assign w6279 = w48499 ^ w48498;
	assign w5569 = w5573 ^ w43765;
	assign w5572 = w43767 ^ w5569;
	assign w5669 = w5571 ^ w5572;
	assign w5568 = w5564 ^ w5569;
	assign w5668 = w5567 ^ w5568;
	assign w43769 = w5774 ^ w5777;
	assign w5687 = w5713 ^ w43769;
	assign w5771 = w5687 ^ w5712;
	assign w5768 = w5769 ^ w5771;
	assign w5727 = w5775 ^ w43769;
	assign w5683 = w5778 ^ w5727;
	assign w5765 = w47803 ^ w5683;
	assign w43772 = w5774 ^ w5780;
	assign w5686 = w5718 ^ w43772;
	assign w5729 = w47799 ^ w5686;
	assign w5764 = w5769 ^ w5729;
	assign w5763 = w5764 & w5765;
	assign w5762 = w5763 ^ w5771;
	assign w5761 = w5769 ^ w5763;
	assign w5682 = w5763 ^ w5727;
	assign w5681 = w5763 ^ w5780;
	assign w5676 = w5681 ^ w5777;
	assign w5760 = w5771 & w5761;
	assign w5758 = w5760 ^ w5768;
	assign w5748 = w5762 & w47804;
	assign w5739 = w5762 & w5794;
	assign w43771 = w5760 ^ w5778;
	assign w5752 = w43771 ^ w5730;
	assign w5750 = w5752 & w5789;
	assign w5741 = w5752 & w5793;
	assign w5719 = w47803 ^ w43771;
	assign w5759 = w5719 ^ w5682;
	assign w5749 = w5759 & w5788;
	assign w5740 = w5759 & w5790;
	assign w5724 = w43772 ^ w5709;
	assign w5770 = w5732 ^ w5724;
	assign w5767 = w5770 & w5768;
	assign w5766 = w5767 ^ w5729;
	assign w5678 = w5767 ^ w5779;
	assign w5674 = w5678 ^ w5714;
	assign w5677 = w47797 ^ w5674;
	assign w5754 = w5676 ^ w5677;
	assign w5675 = w5767 ^ w5723;
	assign w5673 = w47799 ^ w5674;
	assign w5757 = w5766 & w5758;
	assign w5722 = w5757 ^ w5732;
	assign w5756 = w5722 ^ w5724;
	assign w5680 = w5757 ^ w5781;
	assign w5672 = w5719 ^ w5680;
	assign w5679 = w5709 ^ w5672;
	assign w5755 = w5676 ^ w5679;
	assign w5753 = w5722 ^ w5675;
	assign w5751 = w5672 ^ w5673;
	assign w5747 = w5753 & w5783;
	assign w5746 = w5756 & w5795;
	assign w5745 = w5766 & w5785;
	assign w5689 = w5745 ^ w5746;
	assign w5744 = w5754 & w5786;
	assign w5743 = w5751 & w5784;
	assign w5704 = w5743 ^ w5746;
	assign w5701 = ~w5704;
	assign w5700 = w5743 ^ w5744;
	assign w5742 = w5755 & w5787;
	assign w5738 = w5753 & w5798;
	assign w5720 = w5738 ^ w5742;
	assign w5705 = w5747 ^ w5738;
	assign w5698 = ~w5720;
	assign w5737 = w5756 & w5791;
	assign w5707 = w5745 ^ w5737;
	assign w5736 = w5766 & w5792;
	assign w5697 = w5698 ^ w5736;
	assign w5735 = w5754 & w5797;
	assign w5734 = w5751 & w5799;
	assign w5733 = w5755 & w5796;
	assign w5699 = w5744 ^ w5733;
	assign w5695 = ~w5699;
	assign w43770 = w5734 ^ w5735;
	assign w5716 = w5740 ^ w43770;
	assign w5717 = w5741 ^ w5716;
	assign w5721 = w5749 ^ w5717;
	assign w5726 = w5750 ^ w5721;
	assign w5801 = w5726 ^ w5700;
	assign w5690 = w5748 ^ w5721;
	assign w48490 = w5689 ^ w5690;
	assign w5703 = w5707 ^ w43770;
	assign w5702 = w5698 ^ w5703;
	assign w5802 = w5701 ^ w5702;
	assign w43773 = w5746 ^ w5747;
	assign w48491 = w43773 ^ w5726;
	assign w5728 = w5743 ^ w43773;
	assign w5694 = w5739 ^ w5728;
	assign w5691 = ~w5694;
	assign w5688 = w5744 ^ w5728;
	assign w48492 = w5717 ^ w5688;
	assign w43774 = w5748 ^ w5750;
	assign w5706 = w43774 ^ w5703;
	assign w5803 = w5705 ^ w5706;
	assign w5693 = w5697 ^ w43774;
	assign w5696 = w5735 ^ w5693;
	assign w5800 = w5695 ^ w5696;
	assign w5692 = w5716 ^ w5693;
	assign w48489 = w5691 ^ w5692;
	assign w43775 = w5908 ^ w5914;
	assign w5858 = w43775 ^ w5843;
	assign w5904 = w5866 ^ w5858;
	assign w5820 = w5852 ^ w43775;
	assign w5863 = w47783 ^ w5820;
	assign w5898 = w5903 ^ w5863;
	assign w43776 = w5908 ^ w5911;
	assign w5861 = w5909 ^ w43776;
	assign w5817 = w5912 ^ w5861;
	assign w5899 = w47787 ^ w5817;
	assign w5897 = w5898 & w5899;
	assign w5895 = w5903 ^ w5897;
	assign w5816 = w5897 ^ w5861;
	assign w5815 = w5897 ^ w5914;
	assign w5810 = w5815 ^ w5911;
	assign w5821 = w5847 ^ w43776;
	assign w5905 = w5821 ^ w5846;
	assign w5896 = w5897 ^ w5905;
	assign w5902 = w5903 ^ w5905;
	assign w5901 = w5904 & w5902;
	assign w5900 = w5901 ^ w5863;
	assign w5812 = w5901 ^ w5913;
	assign w5808 = w5812 ^ w5848;
	assign w5811 = w47781 ^ w5808;
	assign w5888 = w5810 ^ w5811;
	assign w5809 = w5901 ^ w5857;
	assign w5807 = w47783 ^ w5808;
	assign w5894 = w5905 & w5895;
	assign w5892 = w5894 ^ w5902;
	assign w5891 = w5900 & w5892;
	assign w5856 = w5891 ^ w5866;
	assign w5890 = w5856 ^ w5858;
	assign w5814 = w5891 ^ w5915;
	assign w5887 = w5856 ^ w5809;
	assign w5882 = w5896 & w47788;
	assign w5881 = w5887 & w5917;
	assign w5880 = w5890 & w5929;
	assign w5879 = w5900 & w5919;
	assign w5823 = w5879 ^ w5880;
	assign w5878 = w5888 & w5920;
	assign w5873 = w5896 & w5928;
	assign w5872 = w5887 & w5932;
	assign w5839 = w5881 ^ w5872;
	assign w5871 = w5890 & w5925;
	assign w5841 = w5879 ^ w5871;
	assign w5870 = w5900 & w5926;
	assign w5869 = w5888 & w5931;
	assign w43777 = w5880 ^ w5881;
	assign w43779 = w5894 ^ w5912;
	assign w5853 = w47787 ^ w43779;
	assign w5893 = w5853 ^ w5816;
	assign w5806 = w5853 ^ w5814;
	assign w5813 = w5843 ^ w5806;
	assign w5889 = w5810 ^ w5813;
	assign w5885 = w5806 ^ w5807;
	assign w5883 = w5893 & w5922;
	assign w5877 = w5885 & w5918;
	assign w5838 = w5877 ^ w5880;
	assign w5835 = ~w5838;
	assign w5834 = w5877 ^ w5878;
	assign w5876 = w5889 & w5921;
	assign w5874 = w5893 & w5924;
	assign w5854 = w5872 ^ w5876;
	assign w5832 = ~w5854;
	assign w5831 = w5832 ^ w5870;
	assign w5868 = w5885 & w5933;
	assign w5867 = w5889 & w5930;
	assign w5833 = w5878 ^ w5867;
	assign w5829 = ~w5833;
	assign w43522 = w5868 ^ w5869;
	assign w5850 = w5874 ^ w43522;
	assign w5837 = w5841 ^ w43522;
	assign w5836 = w5832 ^ w5837;
	assign w5936 = w5835 ^ w5836;
	assign w48461 = ~w5936;
	assign w5862 = w5877 ^ w43777;
	assign w5828 = w5873 ^ w5862;
	assign w5825 = ~w5828;
	assign w5822 = w5878 ^ w5862;
	assign w5886 = w43779 ^ w5864;
	assign w5884 = w5886 & w5923;
	assign w5875 = w5886 & w5927;
	assign w5851 = w5875 ^ w5850;
	assign w5855 = w5883 ^ w5851;
	assign w5860 = w5884 ^ w5855;
	assign w48464 = w43777 ^ w5860;
	assign w5935 = w5860 ^ w5834;
	assign w5824 = w5882 ^ w5855;
	assign w48463 = w5823 ^ w5824;
	assign w48465 = w5851 ^ w5822;
	assign w6023 = w48465 ^ w48469;
	assign w6146 = w6161 ^ w48464;
	assign w6258 = ~w6023;
	assign w6271 = ~w48463;
	assign w6259 = w48467 ^ w6271;
	assign w43778 = w5882 ^ w5884;
	assign w5840 = w43778 ^ w5837;
	assign w5937 = w5839 ^ w5840;
	assign w5827 = w5831 ^ w43778;
	assign w5830 = w5869 ^ w5827;
	assign w5934 = w5829 ^ w5830;
	assign w5826 = w5850 ^ w5827;
	assign w48462 = w5825 ^ w5826;
	assign w6261 = w48466 ^ w48462;
	assign w44266 = w21489 ^ w21495;
	assign w21401 = w21433 ^ w44266;
	assign w21444 = w47767 ^ w21401;
	assign w21479 = w21484 ^ w21444;
	assign w21439 = w44266 ^ w21424;
	assign w21485 = w21447 ^ w21439;
	assign w44267 = w21489 ^ w21492;
	assign w21442 = w21490 ^ w44267;
	assign w21398 = w21493 ^ w21442;
	assign w21480 = w47771 ^ w21398;
	assign w21478 = w21479 & w21480;
	assign w21476 = w21484 ^ w21478;
	assign w21396 = w21478 ^ w21495;
	assign w21391 = w21396 ^ w21492;
	assign w21397 = w21478 ^ w21442;
	assign w21402 = w21428 ^ w44267;
	assign w21486 = w21402 ^ w21427;
	assign w21477 = w21478 ^ w21486;
	assign w21483 = w21484 ^ w21486;
	assign w21482 = w21485 & w21483;
	assign w21481 = w21482 ^ w21444;
	assign w21393 = w21482 ^ w21494;
	assign w21389 = w21393 ^ w21429;
	assign w21392 = w47765 ^ w21389;
	assign w21469 = w21391 ^ w21392;
	assign w21390 = w21482 ^ w21438;
	assign w21388 = w47767 ^ w21389;
	assign w21475 = w21486 & w21476;
	assign w21473 = w21475 ^ w21483;
	assign w21472 = w21481 & w21473;
	assign w21437 = w21472 ^ w21447;
	assign w21471 = w21437 ^ w21439;
	assign w21395 = w21472 ^ w21496;
	assign w21468 = w21437 ^ w21390;
	assign w21463 = w21477 & w47772;
	assign w21462 = w21468 & w21498;
	assign w21461 = w21471 & w21510;
	assign w21460 = w21481 & w21500;
	assign w21404 = w21460 ^ w21461;
	assign w21459 = w21469 & w21501;
	assign w21454 = w21477 & w21509;
	assign w21453 = w21468 & w21513;
	assign w21420 = w21462 ^ w21453;
	assign w21452 = w21471 & w21506;
	assign w21422 = w21460 ^ w21452;
	assign w21451 = w21481 & w21507;
	assign w21450 = w21469 & w21512;
	assign w44269 = w21461 ^ w21462;
	assign w44271 = w21475 ^ w21493;
	assign w21467 = w44271 ^ w21445;
	assign w21465 = w21467 & w21504;
	assign w21456 = w21467 & w21508;
	assign w44270 = w21463 ^ w21465;
	assign w21434 = w47771 ^ w44271;
	assign w21474 = w21434 ^ w21397;
	assign w21387 = w21434 ^ w21395;
	assign w21394 = w21424 ^ w21387;
	assign w21470 = w21391 ^ w21394;
	assign w21466 = w21387 ^ w21388;
	assign w21464 = w21474 & w21503;
	assign w21458 = w21466 & w21499;
	assign w21443 = w21458 ^ w44269;
	assign w21419 = w21458 ^ w21461;
	assign w21416 = ~w21419;
	assign w21415 = w21458 ^ w21459;
	assign w21409 = w21454 ^ w21443;
	assign w21406 = ~w21409;
	assign w21403 = w21459 ^ w21443;
	assign w21457 = w21470 & w21502;
	assign w21435 = w21453 ^ w21457;
	assign w21413 = ~w21435;
	assign w21412 = w21413 ^ w21451;
	assign w21408 = w21412 ^ w44270;
	assign w21411 = w21450 ^ w21408;
	assign w21455 = w21474 & w21505;
	assign w21449 = w21466 & w21514;
	assign w21448 = w21470 & w21511;
	assign w21414 = w21459 ^ w21448;
	assign w21410 = ~w21414;
	assign w21515 = w21410 ^ w21411;
	assign w44268 = w21449 ^ w21450;
	assign w21431 = w21455 ^ w44268;
	assign w21432 = w21456 ^ w21431;
	assign w21436 = w21464 ^ w21432;
	assign w21441 = w21465 ^ w21436;
	assign w48508 = w44269 ^ w21441;
	assign w21516 = w21441 ^ w21415;
	assign w21407 = w21431 ^ w21408;
	assign w48506 = w21406 ^ w21407;
	assign w21405 = w21463 ^ w21436;
	assign w48507 = w21404 ^ w21405;
	assign w6265 = w48507 ^ w48506;
	assign w48509 = w21432 ^ w21403;
	assign w21418 = w21422 ^ w44268;
	assign w21421 = w44270 ^ w21418;
	assign w21518 = w21420 ^ w21421;
	assign w21417 = w21413 ^ w21418;
	assign w21517 = w21416 ^ w21417;
	assign w44272 = w21623 ^ w21626;
	assign w21536 = w21562 ^ w44272;
	assign w21620 = w21536 ^ w21561;
	assign w21617 = w21618 ^ w21620;
	assign w21576 = w21624 ^ w44272;
	assign w21532 = w21627 ^ w21576;
	assign w21614 = w47795 ^ w21532;
	assign w44275 = w21623 ^ w21629;
	assign w21535 = w21567 ^ w44275;
	assign w21578 = w47791 ^ w21535;
	assign w21613 = w21618 ^ w21578;
	assign w21612 = w21613 & w21614;
	assign w21611 = w21612 ^ w21620;
	assign w21610 = w21618 ^ w21612;
	assign w21531 = w21612 ^ w21576;
	assign w21530 = w21612 ^ w21629;
	assign w21525 = w21530 ^ w21626;
	assign w21609 = w21620 & w21610;
	assign w21607 = w21609 ^ w21617;
	assign w21597 = w21611 & w47796;
	assign w21588 = w21611 & w21643;
	assign w44274 = w21609 ^ w21627;
	assign w21601 = w44274 ^ w21579;
	assign w21599 = w21601 & w21638;
	assign w21590 = w21601 & w21642;
	assign w21568 = w47795 ^ w44274;
	assign w21608 = w21568 ^ w21531;
	assign w21598 = w21608 & w21637;
	assign w21589 = w21608 & w21639;
	assign w21573 = w44275 ^ w21558;
	assign w21619 = w21581 ^ w21573;
	assign w21616 = w21619 & w21617;
	assign w21615 = w21616 ^ w21578;
	assign w21527 = w21616 ^ w21628;
	assign w21523 = w21527 ^ w21563;
	assign w21526 = w47789 ^ w21523;
	assign w21603 = w21525 ^ w21526;
	assign w21524 = w21616 ^ w21572;
	assign w21522 = w47791 ^ w21523;
	assign w21606 = w21615 & w21607;
	assign w21571 = w21606 ^ w21581;
	assign w21605 = w21571 ^ w21573;
	assign w21529 = w21606 ^ w21630;
	assign w21521 = w21568 ^ w21529;
	assign w21528 = w21558 ^ w21521;
	assign w21604 = w21525 ^ w21528;
	assign w21602 = w21571 ^ w21524;
	assign w21600 = w21521 ^ w21522;
	assign w21596 = w21602 & w21632;
	assign w21595 = w21605 & w21644;
	assign w21594 = w21615 & w21634;
	assign w21538 = w21594 ^ w21595;
	assign w21593 = w21603 & w21635;
	assign w21592 = w21600 & w21633;
	assign w21553 = w21592 ^ w21595;
	assign w21550 = ~w21553;
	assign w21549 = w21592 ^ w21593;
	assign w21591 = w21604 & w21636;
	assign w21587 = w21602 & w21647;
	assign w21569 = w21587 ^ w21591;
	assign w21554 = w21596 ^ w21587;
	assign w21547 = ~w21569;
	assign w21586 = w21605 & w21640;
	assign w21556 = w21594 ^ w21586;
	assign w21585 = w21615 & w21641;
	assign w21546 = w21547 ^ w21585;
	assign w21584 = w21603 & w21646;
	assign w21583 = w21600 & w21648;
	assign w21582 = w21604 & w21645;
	assign w21548 = w21593 ^ w21582;
	assign w21544 = ~w21548;
	assign w44273 = w21583 ^ w21584;
	assign w21565 = w21589 ^ w44273;
	assign w21566 = w21590 ^ w21565;
	assign w21570 = w21598 ^ w21566;
	assign w21575 = w21599 ^ w21570;
	assign w21650 = w21575 ^ w21549;
	assign w21539 = w21597 ^ w21570;
	assign w48475 = w21538 ^ w21539;
	assign w5981 = w48475 ^ w48480;
	assign w6214 = ~w5981;
	assign w6250 = w48481 ^ w48475;
	assign w21552 = w21556 ^ w44273;
	assign w21551 = w21547 ^ w21552;
	assign w21651 = w21550 ^ w21551;
	assign w44276 = w21595 ^ w21596;
	assign w48476 = w44276 ^ w21575;
	assign w5989 = w48476 ^ w48481;
	assign w6173 = w5264 ^ w48476;
	assign w6217 = ~w5989;
	assign w21577 = w21592 ^ w44276;
	assign w21543 = w21588 ^ w21577;
	assign w21540 = ~w21543;
	assign w21537 = w21593 ^ w21577;
	assign w48477 = w21566 ^ w21537;
	assign w6029 = w48477 ^ w48484;
	assign w6024 = w48477 ^ w48492;
	assign w6251 = w6024 ^ w48490;
	assign w5952 = w6251 ^ w6250;
	assign w6255 = ~w6024;
	assign w6254 = w6255 ^ w48489;
	assign w44277 = w21597 ^ w21599;
	assign w21555 = w44277 ^ w21552;
	assign w21652 = w21554 ^ w21555;
	assign w21542 = w21546 ^ w44277;
	assign w21545 = w21584 ^ w21542;
	assign w21649 = w21544 ^ w21545;
	assign w21541 = w21565 ^ w21542;
	assign w48474 = w21540 ^ w21541;
	assign w5974 = w48474 ^ w48479;
	assign w6198 = ~w5974;
	assign w6200 = w6198 ^ w48489;
	assign w6253 = w6252 ^ w48474;
	assign w5951 = w6254 ^ w6253;
	assign w44278 = w21757 ^ w21763;
	assign w21707 = w44278 ^ w21692;
	assign w21753 = w21715 ^ w21707;
	assign w21669 = w21701 ^ w44278;
	assign w21712 = w47807 ^ w21669;
	assign w21747 = w21752 ^ w21712;
	assign w44279 = w21757 ^ w21760;
	assign w21710 = w21758 ^ w44279;
	assign w21666 = w21761 ^ w21710;
	assign w21748 = w47811 ^ w21666;
	assign w21746 = w21747 & w21748;
	assign w21744 = w21752 ^ w21746;
	assign w21665 = w21746 ^ w21710;
	assign w21664 = w21746 ^ w21763;
	assign w21659 = w21664 ^ w21760;
	assign w21670 = w21696 ^ w44279;
	assign w21754 = w21670 ^ w21695;
	assign w21745 = w21746 ^ w21754;
	assign w21751 = w21752 ^ w21754;
	assign w21750 = w21753 & w21751;
	assign w21749 = w21750 ^ w21712;
	assign w21661 = w21750 ^ w21762;
	assign w21657 = w21661 ^ w21697;
	assign w21660 = w47805 ^ w21657;
	assign w21737 = w21659 ^ w21660;
	assign w21658 = w21750 ^ w21706;
	assign w21656 = w47807 ^ w21657;
	assign w21743 = w21754 & w21744;
	assign w21741 = w21743 ^ w21751;
	assign w21740 = w21749 & w21741;
	assign w21705 = w21740 ^ w21715;
	assign w21739 = w21705 ^ w21707;
	assign w21663 = w21740 ^ w21764;
	assign w21736 = w21705 ^ w21658;
	assign w21731 = w21745 & w47812;
	assign w21730 = w21736 & w21766;
	assign w21729 = w21739 & w21778;
	assign w21728 = w21749 & w21768;
	assign w21672 = w21728 ^ w21729;
	assign w21727 = w21737 & w21769;
	assign w21722 = w21745 & w21777;
	assign w21721 = w21736 & w21781;
	assign w21688 = w21730 ^ w21721;
	assign w21720 = w21739 & w21774;
	assign w21690 = w21728 ^ w21720;
	assign w21719 = w21749 & w21775;
	assign w21718 = w21737 & w21780;
	assign w44280 = w21729 ^ w21730;
	assign w44282 = w21743 ^ w21761;
	assign w21702 = w47811 ^ w44282;
	assign w21742 = w21702 ^ w21665;
	assign w21655 = w21702 ^ w21663;
	assign w21662 = w21692 ^ w21655;
	assign w21738 = w21659 ^ w21662;
	assign w21734 = w21655 ^ w21656;
	assign w21732 = w21742 & w21771;
	assign w21726 = w21734 & w21767;
	assign w21687 = w21726 ^ w21729;
	assign w21684 = ~w21687;
	assign w21683 = w21726 ^ w21727;
	assign w21725 = w21738 & w21770;
	assign w21723 = w21742 & w21773;
	assign w21703 = w21721 ^ w21725;
	assign w21681 = ~w21703;
	assign w21680 = w21681 ^ w21719;
	assign w21717 = w21734 & w21782;
	assign w21716 = w21738 & w21779;
	assign w21682 = w21727 ^ w21716;
	assign w21678 = ~w21682;
	assign w43559 = w21717 ^ w21718;
	assign w21699 = w21723 ^ w43559;
	assign w21686 = w21690 ^ w43559;
	assign w21685 = w21681 ^ w21686;
	assign w21785 = w21684 ^ w21685;
	assign w21711 = w21726 ^ w44280;
	assign w21677 = w21722 ^ w21711;
	assign w21674 = ~w21677;
	assign w21671 = w21727 ^ w21711;
	assign w21735 = w44282 ^ w21713;
	assign w21733 = w21735 & w21772;
	assign w21724 = w21735 & w21776;
	assign w21700 = w21724 ^ w21699;
	assign w21704 = w21732 ^ w21700;
	assign w21709 = w21733 ^ w21704;
	assign w48504 = w44280 ^ w21709;
	assign w6017 = w48504 ^ w48508;
	assign w21784 = w21709 ^ w21683;
	assign w21673 = w21731 ^ w21704;
	assign w48503 = w21672 ^ w21673;
	assign w6014 = w48499 ^ w48503;
	assign w6226 = w48504 ^ w48503;
	assign w48505 = w21700 ^ w21671;
	assign w6034 = w48505 ^ w48509;
	assign w6019 = w48501 ^ w48505;
	assign w6062 = w6019 ^ w48508;
	assign w6227 = w6034 ^ w48507;
	assign w5962 = w6227 ^ w6226;
	assign w44281 = w21731 ^ w21733;
	assign w21689 = w44281 ^ w21686;
	assign w21786 = w21688 ^ w21689;
	assign w21676 = w21680 ^ w44281;
	assign w21679 = w21718 ^ w21676;
	assign w21783 = w21678 ^ w21679;
	assign w21675 = w21699 ^ w21676;
	assign w48502 = w21674 ^ w21675;
	assign w6016 = w48502 ^ w48506;
	assign w6075 = w6014 ^ w6016;
	assign w6280 = w6019 ^ w48502;
	assign w5940 = w6280 ^ w6279;
	assign w44283 = w21891 ^ w21897;
	assign w21803 = w21835 ^ w44283;
	assign w21846 = w47839 ^ w21803;
	assign w21881 = w21886 ^ w21846;
	assign w21841 = w44283 ^ w21826;
	assign w21887 = w21849 ^ w21841;
	assign w44284 = w21891 ^ w21894;
	assign w21844 = w21892 ^ w44284;
	assign w21800 = w21895 ^ w21844;
	assign w21882 = w47843 ^ w21800;
	assign w21880 = w21881 & w21882;
	assign w21799 = w21880 ^ w21844;
	assign w21798 = w21880 ^ w21897;
	assign w21793 = w21798 ^ w21894;
	assign w21878 = w21886 ^ w21880;
	assign w21804 = w21830 ^ w44284;
	assign w21888 = w21804 ^ w21829;
	assign w21879 = w21880 ^ w21888;
	assign w21885 = w21886 ^ w21888;
	assign w21884 = w21887 & w21885;
	assign w21883 = w21884 ^ w21846;
	assign w21795 = w21884 ^ w21896;
	assign w21791 = w21795 ^ w21831;
	assign w21794 = w47837 ^ w21791;
	assign w21871 = w21793 ^ w21794;
	assign w21792 = w21884 ^ w21840;
	assign w21790 = w47839 ^ w21791;
	assign w21877 = w21888 & w21878;
	assign w21875 = w21877 ^ w21885;
	assign w21874 = w21883 & w21875;
	assign w21839 = w21874 ^ w21849;
	assign w21873 = w21839 ^ w21841;
	assign w21797 = w21874 ^ w21898;
	assign w21870 = w21839 ^ w21792;
	assign w21865 = w21879 & w47844;
	assign w21864 = w21870 & w21900;
	assign w21863 = w21873 & w21912;
	assign w21862 = w21883 & w21902;
	assign w21806 = w21862 ^ w21863;
	assign w21861 = w21871 & w21903;
	assign w21856 = w21879 & w21911;
	assign w21855 = w21870 & w21915;
	assign w21822 = w21864 ^ w21855;
	assign w21854 = w21873 & w21908;
	assign w21824 = w21862 ^ w21854;
	assign w21853 = w21883 & w21909;
	assign w21852 = w21871 & w21914;
	assign w44286 = w21863 ^ w21864;
	assign w44288 = w21877 ^ w21895;
	assign w21869 = w44288 ^ w21847;
	assign w21867 = w21869 & w21906;
	assign w21858 = w21869 & w21910;
	assign w44287 = w21865 ^ w21867;
	assign w21836 = w47843 ^ w44288;
	assign w21876 = w21836 ^ w21799;
	assign w21789 = w21836 ^ w21797;
	assign w21796 = w21826 ^ w21789;
	assign w21872 = w21793 ^ w21796;
	assign w21868 = w21789 ^ w21790;
	assign w21866 = w21876 & w21905;
	assign w21860 = w21868 & w21901;
	assign w21845 = w21860 ^ w44286;
	assign w21821 = w21860 ^ w21863;
	assign w21818 = ~w21821;
	assign w21817 = w21860 ^ w21861;
	assign w21811 = w21856 ^ w21845;
	assign w21808 = ~w21811;
	assign w21805 = w21861 ^ w21845;
	assign w21859 = w21872 & w21904;
	assign w21837 = w21855 ^ w21859;
	assign w21815 = ~w21837;
	assign w21814 = w21815 ^ w21853;
	assign w21810 = w21814 ^ w44287;
	assign w21813 = w21852 ^ w21810;
	assign w21857 = w21876 & w21907;
	assign w21851 = w21868 & w21916;
	assign w21850 = w21872 & w21913;
	assign w21816 = w21861 ^ w21850;
	assign w21812 = ~w21816;
	assign w21917 = w21812 ^ w21813;
	assign w44285 = w21851 ^ w21852;
	assign w21833 = w21857 ^ w44285;
	assign w21834 = w21858 ^ w21833;
	assign w21838 = w21866 ^ w21834;
	assign w21843 = w21867 ^ w21838;
	assign w48487 = w44286 ^ w21843;
	assign w6001 = w48487 ^ w48491;
	assign w48377 = w5952 ^ w6001;
	assign w47696 = w48377 ^ w68;
	assign w6191 = w6214 ^ w6001;
	assign w6201 = w48487 ^ w48481;
	assign w21918 = w21843 ^ w21817;
	assign w21809 = w21833 ^ w21810;
	assign w48485 = w21808 ^ w21809;
	assign w5982 = w48485 ^ w48489;
	assign w6169 = ~w5982;
	assign w6216 = w6214 ^ w5982;
	assign w6246 = w48485 ^ w6245;
	assign w21807 = w21865 ^ w21838;
	assign w48486 = w21806 ^ w21807;
	assign w5992 = w48486 ^ w48490;
	assign w48376 = w5951 ^ w5992;
	assign w47697 = w48376 ^ w67;
	assign w6189 = w6198 ^ w5992;
	assign w6219 = w6217 ^ w5992;
	assign w6242 = w48486 ^ w6252;
	assign w48488 = w21834 ^ w21805;
	assign w6032 = w48488 ^ w48492;
	assign w6025 = w48484 ^ w48488;
	assign w6244 = ~w6025;
	assign w6243 = w6244 ^ w48491;
	assign w5955 = w6243 ^ w6242;
	assign w48393 = w5955 ^ w5989;
	assign w47680 = w48393 ^ w84;
	assign w6247 = w6244 ^ w48490;
	assign w5954 = w6247 ^ w6246;
	assign w48392 = w5954 ^ w5981;
	assign w47681 = w48392 ^ w83;
	assign w21820 = w21824 ^ w44285;
	assign w21823 = w44287 ^ w21820;
	assign w21920 = w21822 ^ w21823;
	assign w21819 = w21815 ^ w21820;
	assign w21919 = w21818 ^ w21819;
	assign w44289 = w22025 ^ w22028;
	assign w21938 = w21964 ^ w44289;
	assign w22022 = w21938 ^ w21963;
	assign w22019 = w22020 ^ w22022;
	assign w21978 = w22026 ^ w44289;
	assign w21934 = w22029 ^ w21978;
	assign w22016 = w47859 ^ w21934;
	assign w44292 = w22025 ^ w22031;
	assign w21937 = w21969 ^ w44292;
	assign w21980 = w47855 ^ w21937;
	assign w22015 = w22020 ^ w21980;
	assign w22014 = w22015 & w22016;
	assign w22013 = w22014 ^ w22022;
	assign w22012 = w22020 ^ w22014;
	assign w21933 = w22014 ^ w21978;
	assign w21932 = w22014 ^ w22031;
	assign w21927 = w21932 ^ w22028;
	assign w22011 = w22022 & w22012;
	assign w22009 = w22011 ^ w22019;
	assign w21999 = w22013 & w47860;
	assign w21990 = w22013 & w22045;
	assign w44291 = w22011 ^ w22029;
	assign w22003 = w44291 ^ w21981;
	assign w22001 = w22003 & w22040;
	assign w21992 = w22003 & w22044;
	assign w21970 = w47859 ^ w44291;
	assign w22010 = w21970 ^ w21933;
	assign w22000 = w22010 & w22039;
	assign w21991 = w22010 & w22041;
	assign w21975 = w44292 ^ w21960;
	assign w22021 = w21983 ^ w21975;
	assign w22018 = w22021 & w22019;
	assign w22017 = w22018 ^ w21980;
	assign w21929 = w22018 ^ w22030;
	assign w21925 = w21929 ^ w21965;
	assign w21928 = w47853 ^ w21925;
	assign w22005 = w21927 ^ w21928;
	assign w21926 = w22018 ^ w21974;
	assign w21924 = w47855 ^ w21925;
	assign w22008 = w22017 & w22009;
	assign w21973 = w22008 ^ w21983;
	assign w22007 = w21973 ^ w21975;
	assign w21931 = w22008 ^ w22032;
	assign w21923 = w21970 ^ w21931;
	assign w21930 = w21960 ^ w21923;
	assign w22006 = w21927 ^ w21930;
	assign w22004 = w21973 ^ w21926;
	assign w22002 = w21923 ^ w21924;
	assign w21998 = w22004 & w22034;
	assign w21997 = w22007 & w22046;
	assign w21996 = w22017 & w22036;
	assign w21940 = w21996 ^ w21997;
	assign w21995 = w22005 & w22037;
	assign w21994 = w22002 & w22035;
	assign w21955 = w21994 ^ w21997;
	assign w21952 = ~w21955;
	assign w21951 = w21994 ^ w21995;
	assign w21993 = w22006 & w22038;
	assign w21989 = w22004 & w22049;
	assign w21971 = w21989 ^ w21993;
	assign w21956 = w21998 ^ w21989;
	assign w21949 = ~w21971;
	assign w21988 = w22007 & w22042;
	assign w21958 = w21996 ^ w21988;
	assign w21987 = w22017 & w22043;
	assign w21948 = w21949 ^ w21987;
	assign w21986 = w22005 & w22048;
	assign w21985 = w22002 & w22050;
	assign w21984 = w22006 & w22047;
	assign w21950 = w21995 ^ w21984;
	assign w21946 = ~w21950;
	assign w44290 = w21985 ^ w21986;
	assign w21967 = w21991 ^ w44290;
	assign w21968 = w21992 ^ w21967;
	assign w21972 = w22000 ^ w21968;
	assign w21977 = w22001 ^ w21972;
	assign w22052 = w21977 ^ w21951;
	assign w21941 = w21999 ^ w21972;
	assign w48438 = w21940 ^ w21941;
	assign w21954 = w21958 ^ w44290;
	assign w21953 = w21949 ^ w21954;
	assign w22053 = w21952 ^ w21953;
	assign w44293 = w21997 ^ w21998;
	assign w48439 = w44293 ^ w21977;
	assign w21979 = w21994 ^ w44293;
	assign w21945 = w21990 ^ w21979;
	assign w21942 = ~w21945;
	assign w21939 = w21995 ^ w21979;
	assign w48440 = w21968 ^ w21939;
	assign w6020 = w48440 ^ w48456;
	assign w6124 = ~w6020;
	assign w6278 = w6020 ^ w48438;
	assign w44294 = w21999 ^ w22001;
	assign w21957 = w44294 ^ w21954;
	assign w22054 = w21956 ^ w21957;
	assign w21944 = w21948 ^ w44294;
	assign w21947 = w21986 ^ w21944;
	assign w22051 = w21946 ^ w21947;
	assign w21943 = w21967 ^ w21944;
	assign w48437 = w21942 ^ w21943;
	assign w5985 = w48437 ^ w48452;
	assign w6123 = ~w5985;
	assign w44346 = w23365 ^ w23371;
	assign w23315 = w44346 ^ w23300;
	assign w23361 = w23323 ^ w23315;
	assign w23277 = w23309 ^ w44346;
	assign w23320 = w1442 ^ w23277;
	assign w23355 = w23360 ^ w23320;
	assign w44347 = w23365 ^ w23368;
	assign w23318 = w23366 ^ w44347;
	assign w23274 = w23369 ^ w23318;
	assign w23356 = w1438 ^ w23274;
	assign w23354 = w23355 & w23356;
	assign w23352 = w23360 ^ w23354;
	assign w23273 = w23354 ^ w23318;
	assign w23272 = w23354 ^ w23371;
	assign w23267 = w23272 ^ w23368;
	assign w23278 = w23304 ^ w44347;
	assign w23362 = w23278 ^ w23303;
	assign w23353 = w23354 ^ w23362;
	assign w23359 = w23360 ^ w23362;
	assign w23358 = w23361 & w23359;
	assign w23357 = w23358 ^ w23320;
	assign w23269 = w23358 ^ w23370;
	assign w23265 = w23269 ^ w23305;
	assign w23268 = w1444 ^ w23265;
	assign w23345 = w23267 ^ w23268;
	assign w23266 = w23358 ^ w23314;
	assign w23264 = w1442 ^ w23265;
	assign w23351 = w23362 & w23352;
	assign w23349 = w23351 ^ w23359;
	assign w23348 = w23357 & w23349;
	assign w23313 = w23348 ^ w23323;
	assign w23347 = w23313 ^ w23315;
	assign w23271 = w23348 ^ w23372;
	assign w23344 = w23313 ^ w23266;
	assign w23339 = w23353 & w1437;
	assign w23338 = w23344 & w23374;
	assign w23337 = w23347 & w23386;
	assign w23336 = w23357 & w23376;
	assign w23280 = w23336 ^ w23337;
	assign w23335 = w23345 & w23377;
	assign w23330 = w23353 & w23385;
	assign w23329 = w23344 & w23389;
	assign w23296 = w23338 ^ w23329;
	assign w23328 = w23347 & w23382;
	assign w23298 = w23336 ^ w23328;
	assign w23327 = w23357 & w23383;
	assign w23326 = w23345 & w23388;
	assign w44348 = w23337 ^ w23338;
	assign w44350 = w23351 ^ w23369;
	assign w23310 = w1438 ^ w44350;
	assign w23350 = w23310 ^ w23273;
	assign w23263 = w23310 ^ w23271;
	assign w23270 = w23300 ^ w23263;
	assign w23346 = w23267 ^ w23270;
	assign w23342 = w23263 ^ w23264;
	assign w23340 = w23350 & w23379;
	assign w23334 = w23342 & w23375;
	assign w23295 = w23334 ^ w23337;
	assign w23292 = ~w23295;
	assign w23291 = w23334 ^ w23335;
	assign w23333 = w23346 & w23378;
	assign w23331 = w23350 & w23381;
	assign w23311 = w23329 ^ w23333;
	assign w23289 = ~w23311;
	assign w23288 = w23289 ^ w23327;
	assign w23325 = w23342 & w23390;
	assign w23324 = w23346 & w23387;
	assign w23290 = w23335 ^ w23324;
	assign w23286 = ~w23290;
	assign w43563 = w23325 ^ w23326;
	assign w23307 = w23331 ^ w43563;
	assign w23294 = w23298 ^ w43563;
	assign w23293 = w23289 ^ w23294;
	assign w23393 = w23292 ^ w23293;
	assign w47966 = ~w23393;
	assign w1478 = w1892 ^ w47966;
	assign w1509 = w1923 ^ w1478;
	assign w1541 = w1955 ^ w1509;
	assign w1573 = w1987 ^ w1541;
	assign w23319 = w23334 ^ w44348;
	assign w23285 = w23330 ^ w23319;
	assign w23282 = ~w23285;
	assign w23279 = w23335 ^ w23319;
	assign w23343 = w44350 ^ w23321;
	assign w23341 = w23343 & w23380;
	assign w23332 = w23343 & w23384;
	assign w23308 = w23332 ^ w23307;
	assign w23312 = w23340 ^ w23308;
	assign w23317 = w23341 ^ w23312;
	assign w47969 = w44348 ^ w23317;
	assign w1481 = w1895 ^ w47969;
	assign w1512 = w1926 ^ w1481;
	assign w1544 = w1958 ^ w1512;
	assign w1576 = w1990 ^ w1544;
	assign w23392 = w23317 ^ w23291;
	assign w23281 = w23339 ^ w23312;
	assign w47968 = w23280 ^ w23281;
	assign w1480 = w1894 ^ w47968;
	assign w1511 = w1925 ^ w1480;
	assign w1543 = w1957 ^ w1511;
	assign w1575 = w1989 ^ w1543;
	assign w4768 = w1573 ^ w1575;
	assign w47972 = w23308 ^ w23279;
	assign w1484 = w1898 ^ w47972;
	assign w1515 = w1929 ^ w1484;
	assign w1547 = w1961 ^ w1515;
	assign w1579 = w1993 ^ w1547;
	assign w4858 = w1576 ^ w1579;
	assign w4850 = w4768 ^ w4858;
	assign w4859 = w1579 ^ w1573;
	assign w47971 = ~w23392;
	assign w1483 = w1897 ^ w47971;
	assign w1514 = w1928 ^ w1483;
	assign w1546 = w1960 ^ w1514;
	assign w1578 = w1992 ^ w1546;
	assign w4771 = w1576 ^ w1578;
	assign w44349 = w23339 ^ w23341;
	assign w23297 = w44349 ^ w23294;
	assign w23394 = w23296 ^ w23297;
	assign w47965 = ~w23394;
	assign w1477 = w1891 ^ w47965;
	assign w1508 = w1922 ^ w1477;
	assign w1540 = w1954 ^ w1508;
	assign w1572 = w1986 ^ w1540;
	assign w4849 = w1572 ^ w4850;
	assign w4775 = w1572 ^ w1578;
	assign w23284 = w23288 ^ w44349;
	assign w23287 = w23326 ^ w23284;
	assign w23391 = w23286 ^ w23287;
	assign w23283 = w23307 ^ w23284;
	assign w47967 = w23282 ^ w23283;
	assign w1479 = w1893 ^ w47967;
	assign w1510 = w1924 ^ w1479;
	assign w1542 = w1956 ^ w1510;
	assign w1574 = w1988 ^ w1542;
	assign w4770 = w1574 ^ w4768;
	assign w4847 = w1578 ^ w4770;
	assign w4846 = w4775 ^ w4770;
	assign w4785 = w1573 ^ w1574;
	assign w4854 = w4858 ^ w4785;
	assign w4860 = w1574 ^ w1576;
	assign w4745 = w1575 ^ w1574;
	assign w4857 = w1579 ^ w1574;
	assign w4843 = w4850 & w4854;
	assign w4774 = w4843 ^ w4771;
	assign w4837 = w4858 & w4847;
	assign w4772 = w4837 ^ w4770;
	assign w4778 = w4774 ^ w4772;
	assign w4783 = w1579 ^ w4778;
	assign w47970 = ~w23391;
	assign w1482 = w1896 ^ w47970;
	assign w1513 = w1927 ^ w1482;
	assign w1545 = w1959 ^ w1513;
	assign w1577 = w1991 ^ w1545;
	assign w4844 = w1577 ^ w4770;
	assign w4769 = w1577 ^ w1579;
	assign w4845 = w4769 ^ w4860;
	assign w4853 = w4769 ^ w4775;
	assign w4851 = w4785 ^ w4853;
	assign w4856 = w1577 ^ w4775;
	assign w4852 = w1573 ^ w4856;
	assign w4731 = w4771 ^ w4769;
	assign w4848 = w4768 ^ w4731;
	assign w4730 = w4771 ^ w1577;
	assign w4855 = w1572 ^ w4730;
	assign w4842 = w4851 & w4849;
	assign w4841 = w4855 & w1572;
	assign w4840 = w4859 & w4844;
	assign w4773 = w4840 ^ w4769;
	assign w4839 = w4856 & w4852;
	assign w4838 = w4853 & w4846;
	assign w4836 = w4860 & w4845;
	assign w4792 = w4836 ^ w4842;
	assign w4834 = w4792 ^ w4783;
	assign w4744 = w4836 ^ w4837;
	assign w4791 = w4744 ^ w4745;
	assign w4790 = w4791 ^ w4773;
	assign w4833 = w4839 ^ w4790;
	assign w4835 = w4857 & w4848;
	assign w4830 = w4834 & w4833;
	assign w43519 = w4835 ^ w4838;
	assign w4787 = w4836 ^ w43519;
	assign w4743 = w4839 ^ w4787;
	assign w4826 = w1573 ^ w4743;
	assign w4747 = w4773 ^ w43519;
	assign w4832 = w4747 ^ w4772;
	assign w4829 = w4830 ^ w4832;
	assign w43733 = w4835 ^ w4841;
	assign w4746 = w4778 ^ w43733;
	assign w4789 = w1577 ^ w4746;
	assign w4825 = w4830 ^ w4789;
	assign w4824 = w4825 & w4826;
	assign w4822 = w4830 ^ w4824;
	assign w4742 = w4824 ^ w4787;
	assign w4741 = w4824 ^ w4841;
	assign w4736 = w4741 ^ w4838;
	assign w4823 = w4824 ^ w4832;
	assign w4821 = w4832 & w4822;
	assign w4819 = w4821 ^ w4829;
	assign w4809 = w4823 & w1572;
	assign w4800 = w4823 & w4855;
	assign w43732 = w4821 ^ w4839;
	assign w4813 = w43732 ^ w4790;
	assign w4811 = w4813 & w4850;
	assign w4802 = w4813 & w4854;
	assign w4779 = w1573 ^ w43732;
	assign w4820 = w4779 ^ w4742;
	assign w4810 = w4820 & w4849;
	assign w4801 = w4820 & w4851;
	assign w4784 = w43733 ^ w4769;
	assign w4831 = w4792 ^ w4784;
	assign w4828 = w4831 & w4829;
	assign w4827 = w4828 ^ w4789;
	assign w4738 = w4828 ^ w4840;
	assign w4734 = w4738 ^ w4774;
	assign w4737 = w1579 ^ w4734;
	assign w4815 = w4736 ^ w4737;
	assign w4735 = w4828 ^ w4783;
	assign w4733 = w1577 ^ w4734;
	assign w4818 = w4827 & w4819;
	assign w4782 = w4818 ^ w4792;
	assign w4817 = w4782 ^ w4784;
	assign w4740 = w4818 ^ w4842;
	assign w4732 = w4779 ^ w4740;
	assign w4739 = w4769 ^ w4732;
	assign w4816 = w4736 ^ w4739;
	assign w4814 = w4782 ^ w4735;
	assign w4812 = w4732 ^ w4733;
	assign w4808 = w4814 & w4844;
	assign w4807 = w4817 & w4856;
	assign w4806 = w4827 & w4846;
	assign w4749 = w4806 ^ w4807;
	assign w4805 = w4815 & w4847;
	assign w4804 = w4812 & w4845;
	assign w4764 = w4804 ^ w4807;
	assign w4761 = ~w4764;
	assign w4760 = w4804 ^ w4805;
	assign w4803 = w4816 & w4848;
	assign w4799 = w4814 & w4859;
	assign w4780 = w4799 ^ w4803;
	assign w4765 = w4808 ^ w4799;
	assign w4758 = ~w4780;
	assign w4798 = w4817 & w4852;
	assign w4767 = w4806 ^ w4798;
	assign w4797 = w4827 & w4853;
	assign w4757 = w4758 ^ w4797;
	assign w4796 = w4815 & w4858;
	assign w4795 = w4812 & w4860;
	assign w4793 = w4795 ^ w4796;
	assign w4776 = w4801 ^ w4793;
	assign w4777 = w4802 ^ w4776;
	assign w4781 = w4810 ^ w4777;
	assign w4786 = w4811 ^ w4781;
	assign w4763 = w4767 ^ w4793;
	assign w4762 = w4758 ^ w4763;
	assign w4863 = w4761 ^ w4762;
	assign w4862 = w4786 ^ w4760;
	assign w4750 = w4809 ^ w4781;
	assign w48000 = w4749 ^ w4750;
	assign w4794 = w4816 & w4857;
	assign w4759 = w4805 ^ w4794;
	assign w4755 = ~w4759;
	assign w47998 = ~w4863;
	assign w48003 = ~w4862;
	assign w1605 = w2019 ^ w47998;
	assign w1637 = w1382 ^ w1605;
	assign w1610 = w2024 ^ w48003;
	assign w1642 = w1387 ^ w1610;
	assign w1607 = w2021 ^ w48000;
	assign w1639 = w1384 ^ w1607;
	assign w1674 = w1419 ^ w1642;
	assign w1706 = w1451 ^ w1674;
	assign w1671 = w1416 ^ w1639;
	assign w1703 = w1448 ^ w1671;
	assign w1669 = w1414 ^ w1637;
	assign w1701 = w1446 ^ w1669;
	assign w35493 = w1701 ^ w1703;
	assign w43734 = w4807 ^ w4808;
	assign w48001 = w43734 ^ w4786;
	assign w1608 = w2022 ^ w48001;
	assign w1640 = w1385 ^ w1608;
	assign w1672 = w1417 ^ w1640;
	assign w1704 = w1449 ^ w1672;
	assign w35496 = w1704 ^ w1706;
	assign w4788 = w4804 ^ w43734;
	assign w4754 = w4800 ^ w4788;
	assign w4751 = ~w4754;
	assign w4748 = w4805 ^ w4788;
	assign w48004 = w4777 ^ w4748;
	assign w1611 = w2025 ^ w48004;
	assign w1643 = w1388 ^ w1611;
	assign w1675 = w1420 ^ w1643;
	assign w1707 = w1452 ^ w1675;
	assign w35582 = w1704 ^ w1707;
	assign w35574 = w35493 ^ w35582;
	assign w35583 = w1707 ^ w1701;
	assign w43735 = w4809 ^ w4811;
	assign w4753 = w4757 ^ w43735;
	assign w4752 = w4776 ^ w4753;
	assign w4756 = w4796 ^ w4753;
	assign w4861 = w4755 ^ w4756;
	assign w48002 = ~w4861;
	assign w1609 = w2023 ^ w48002;
	assign w1641 = w1386 ^ w1609;
	assign w1673 = w1418 ^ w1641;
	assign w1705 = w1450 ^ w1673;
	assign w35455 = w35496 ^ w1705;
	assign w47999 = w4751 ^ w4752;
	assign w1606 = w2020 ^ w47999;
	assign w1638 = w1383 ^ w1606;
	assign w1670 = w1415 ^ w1638;
	assign w1702 = w1447 ^ w1670;
	assign w35494 = w1705 ^ w1707;
	assign w35495 = w1702 ^ w35493;
	assign w35571 = w1706 ^ w35495;
	assign w35568 = w1705 ^ w35495;
	assign w35510 = w1701 ^ w1702;
	assign w35578 = w35582 ^ w35510;
	assign w35584 = w1702 ^ w1704;
	assign w35569 = w35494 ^ w35584;
	assign w35470 = w1703 ^ w1702;
	assign w35456 = w35496 ^ w35494;
	assign w35572 = w35493 ^ w35456;
	assign w35581 = w1707 ^ w1702;
	assign w35567 = w35574 & w35578;
	assign w35499 = w35567 ^ w35496;
	assign w35564 = w35583 & w35568;
	assign w35498 = w35564 ^ w35494;
	assign w35561 = w35582 & w35571;
	assign w35497 = w35561 ^ w35495;
	assign w35503 = w35499 ^ w35497;
	assign w35508 = w1707 ^ w35503;
	assign w35560 = w35584 & w35569;
	assign w35469 = w35560 ^ w35561;
	assign w35516 = w35469 ^ w35470;
	assign w35515 = w35516 ^ w35498;
	assign w35559 = w35581 & w35572;
	assign w4766 = w43735 ^ w4763;
	assign w4864 = w4765 ^ w4766;
	assign w47997 = ~w4864;
	assign w1604 = w2018 ^ w47997;
	assign w1636 = w1381 ^ w1604;
	assign w1668 = w1413 ^ w1636;
	assign w1700 = w1445 ^ w1668;
	assign w35573 = w1700 ^ w35574;
	assign w35500 = w1700 ^ w1706;
	assign w35570 = w35500 ^ w35495;
	assign w35577 = w35494 ^ w35500;
	assign w35575 = w35510 ^ w35577;
	assign w35580 = w1705 ^ w35500;
	assign w35576 = w1701 ^ w35580;
	assign w35579 = w1700 ^ w35455;
	assign w35566 = w35575 & w35573;
	assign w35517 = w35560 ^ w35566;
	assign w35558 = w35517 ^ w35508;
	assign w35565 = w35579 & w1700;
	assign w35563 = w35580 & w35576;
	assign w35557 = w35563 ^ w35515;
	assign w35562 = w35577 & w35570;
	assign w35554 = w35558 & w35557;
	assign w44452 = w25911 ^ w25917;
	assign w25861 = w44452 ^ w25846;
	assign w25907 = w25869 ^ w25861;
	assign w25823 = w25855 ^ w44452;
	assign w25866 = w47823 ^ w25823;
	assign w25901 = w25906 ^ w25866;
	assign w44453 = w25911 ^ w25914;
	assign w25864 = w25912 ^ w44453;
	assign w25820 = w25915 ^ w25864;
	assign w25902 = w47827 ^ w25820;
	assign w25900 = w25901 & w25902;
	assign w25898 = w25906 ^ w25900;
	assign w25819 = w25900 ^ w25864;
	assign w25818 = w25900 ^ w25917;
	assign w25813 = w25818 ^ w25914;
	assign w25824 = w25850 ^ w44453;
	assign w25908 = w25824 ^ w25849;
	assign w25899 = w25900 ^ w25908;
	assign w25905 = w25906 ^ w25908;
	assign w25904 = w25907 & w25905;
	assign w25903 = w25904 ^ w25866;
	assign w25815 = w25904 ^ w25916;
	assign w25811 = w25815 ^ w25851;
	assign w25814 = w47821 ^ w25811;
	assign w25891 = w25813 ^ w25814;
	assign w25812 = w25904 ^ w25860;
	assign w25810 = w47823 ^ w25811;
	assign w25897 = w25908 & w25898;
	assign w25895 = w25897 ^ w25905;
	assign w25894 = w25903 & w25895;
	assign w25859 = w25894 ^ w25869;
	assign w25893 = w25859 ^ w25861;
	assign w25817 = w25894 ^ w25918;
	assign w25890 = w25859 ^ w25812;
	assign w25885 = w25899 & w47828;
	assign w25884 = w25890 & w25920;
	assign w25883 = w25893 & w25932;
	assign w25882 = w25903 & w25922;
	assign w25826 = w25882 ^ w25883;
	assign w25881 = w25891 & w25923;
	assign w25876 = w25899 & w25931;
	assign w25875 = w25890 & w25935;
	assign w25842 = w25884 ^ w25875;
	assign w25874 = w25893 & w25928;
	assign w25844 = w25882 ^ w25874;
	assign w25873 = w25903 & w25929;
	assign w25872 = w25891 & w25934;
	assign w44454 = w25883 ^ w25884;
	assign w44456 = w25897 ^ w25915;
	assign w25856 = w47827 ^ w44456;
	assign w25896 = w25856 ^ w25819;
	assign w25809 = w25856 ^ w25817;
	assign w25816 = w25846 ^ w25809;
	assign w25892 = w25813 ^ w25816;
	assign w25888 = w25809 ^ w25810;
	assign w25886 = w25896 & w25925;
	assign w25880 = w25888 & w25921;
	assign w25865 = w25880 ^ w44454;
	assign w25841 = w25880 ^ w25883;
	assign w25838 = ~w25841;
	assign w25837 = w25880 ^ w25881;
	assign w25825 = w25881 ^ w25865;
	assign w25879 = w25892 & w25924;
	assign w25877 = w25896 & w25927;
	assign w25831 = w25876 ^ w25865;
	assign w25828 = ~w25831;
	assign w25857 = w25875 ^ w25879;
	assign w25835 = ~w25857;
	assign w25834 = w25835 ^ w25873;
	assign w25871 = w25888 & w25936;
	assign w25870 = w25892 & w25933;
	assign w25836 = w25881 ^ w25870;
	assign w25832 = ~w25836;
	assign w43571 = w25871 ^ w25872;
	assign w25840 = w25844 ^ w43571;
	assign w25839 = w25835 ^ w25840;
	assign w25939 = w25838 ^ w25839;
	assign w25853 = w25877 ^ w43571;
	assign w25889 = w44456 ^ w25867;
	assign w25887 = w25889 & w25926;
	assign w25878 = w25889 & w25930;
	assign w25854 = w25878 ^ w25853;
	assign w25858 = w25886 ^ w25854;
	assign w25863 = w25887 ^ w25858;
	assign w48459 = w44454 ^ w25863;
	assign w6002 = w48459 ^ w48464;
	assign w6160 = ~w6002;
	assign w25938 = w25863 ^ w25837;
	assign w25827 = w25885 ^ w25858;
	assign w48458 = w25826 ^ w25827;
	assign w5998 = w48458 ^ w48463;
	assign w6134 = ~w5998;
	assign w6269 = w48464 ^ w48458;
	assign w48460 = w25854 ^ w25825;
	assign w6030 = w48460 ^ w48465;
	assign w44455 = w25885 ^ w25887;
	assign w25843 = w44455 ^ w25840;
	assign w25940 = w25842 ^ w25843;
	assign w25830 = w25834 ^ w44455;
	assign w25833 = w25872 ^ w25830;
	assign w25937 = w25832 ^ w25833;
	assign w25829 = w25853 ^ w25830;
	assign w48457 = w25828 ^ w25829;
	assign w5995 = w48457 ^ w48462;
	assign w6142 = ~w5995;
	assign w6272 = w6271 ^ w48457;
	assign w44580 = w28993 ^ w28996;
	assign w28906 = w28932 ^ w44580;
	assign w28990 = w28906 ^ w28931;
	assign w28987 = w28988 ^ w28990;
	assign w28946 = w28994 ^ w44580;
	assign w28902 = w28997 ^ w28946;
	assign w28984 = w47779 ^ w28902;
	assign w44583 = w28993 ^ w28999;
	assign w28905 = w28937 ^ w44583;
	assign w28948 = w47775 ^ w28905;
	assign w28983 = w28988 ^ w28948;
	assign w28982 = w28983 & w28984;
	assign w28981 = w28982 ^ w28990;
	assign w28980 = w28988 ^ w28982;
	assign w28901 = w28982 ^ w28946;
	assign w28900 = w28982 ^ w28999;
	assign w28895 = w28900 ^ w28996;
	assign w28979 = w28990 & w28980;
	assign w28977 = w28979 ^ w28987;
	assign w28967 = w28981 & w47780;
	assign w28958 = w28981 & w29013;
	assign w44582 = w28979 ^ w28997;
	assign w28971 = w44582 ^ w28949;
	assign w28969 = w28971 & w29008;
	assign w28960 = w28971 & w29012;
	assign w28938 = w47779 ^ w44582;
	assign w28978 = w28938 ^ w28901;
	assign w28968 = w28978 & w29007;
	assign w28959 = w28978 & w29009;
	assign w28943 = w44583 ^ w28928;
	assign w28989 = w28951 ^ w28943;
	assign w28986 = w28989 & w28987;
	assign w28985 = w28986 ^ w28948;
	assign w28897 = w28986 ^ w28998;
	assign w28893 = w28897 ^ w28933;
	assign w28896 = w47773 ^ w28893;
	assign w28973 = w28895 ^ w28896;
	assign w28894 = w28986 ^ w28942;
	assign w28892 = w47775 ^ w28893;
	assign w28976 = w28985 & w28977;
	assign w28941 = w28976 ^ w28951;
	assign w28975 = w28941 ^ w28943;
	assign w28899 = w28976 ^ w29000;
	assign w28891 = w28938 ^ w28899;
	assign w28898 = w28928 ^ w28891;
	assign w28974 = w28895 ^ w28898;
	assign w28972 = w28941 ^ w28894;
	assign w28970 = w28891 ^ w28892;
	assign w28966 = w28972 & w29002;
	assign w28965 = w28975 & w29014;
	assign w28964 = w28985 & w29004;
	assign w28908 = w28964 ^ w28965;
	assign w28963 = w28973 & w29005;
	assign w28962 = w28970 & w29003;
	assign w28923 = w28962 ^ w28965;
	assign w28920 = ~w28923;
	assign w28919 = w28962 ^ w28963;
	assign w28961 = w28974 & w29006;
	assign w28957 = w28972 & w29017;
	assign w28939 = w28957 ^ w28961;
	assign w28924 = w28966 ^ w28957;
	assign w28917 = ~w28939;
	assign w28956 = w28975 & w29010;
	assign w28926 = w28964 ^ w28956;
	assign w28955 = w28985 & w29011;
	assign w28916 = w28917 ^ w28955;
	assign w28954 = w28973 & w29016;
	assign w28953 = w28970 & w29018;
	assign w28952 = w28974 & w29015;
	assign w28918 = w28963 ^ w28952;
	assign w28914 = ~w28918;
	assign w44581 = w28953 ^ w28954;
	assign w28935 = w28959 ^ w44581;
	assign w28936 = w28960 ^ w28935;
	assign w28940 = w28968 ^ w28936;
	assign w28945 = w28969 ^ w28940;
	assign w29020 = w28945 ^ w28919;
	assign w28909 = w28967 ^ w28940;
	assign w48449 = w28908 ^ w28909;
	assign w5973 = w48449 ^ w48453;
	assign w6126 = w5973 ^ w6123;
	assign w28922 = w28926 ^ w44581;
	assign w28921 = w28917 ^ w28922;
	assign w29021 = w28920 ^ w28921;
	assign w48447 = ~w29021;
	assign w44584 = w28965 ^ w28966;
	assign w48450 = w44584 ^ w28945;
	assign w5976 = w48450 ^ w48454;
	assign w28947 = w28962 ^ w44584;
	assign w28913 = w28958 ^ w28947;
	assign w28910 = ~w28913;
	assign w28907 = w28963 ^ w28947;
	assign w48451 = w28936 ^ w28907;
	assign w6028 = w48451 ^ w48456;
	assign w44585 = w28967 ^ w28969;
	assign w28925 = w44585 ^ w28922;
	assign w29022 = w28924 ^ w28925;
	assign w28912 = w28916 ^ w44585;
	assign w28915 = w28954 ^ w28912;
	assign w29019 = w28914 ^ w28915;
	assign w28911 = w28935 ^ w28912;
	assign w48448 = w28910 ^ w28911;
	assign w6231 = ~w48448;
	assign w6232 = w48449 ^ w6231;
	assign w44733 = w32611 ^ w32617;
	assign w32561 = w44733 ^ w32546;
	assign w32607 = w32569 ^ w32561;
	assign w32523 = w32555 ^ w44733;
	assign w32566 = w47831 ^ w32523;
	assign w32601 = w32606 ^ w32566;
	assign w44734 = w32611 ^ w32614;
	assign w32564 = w32612 ^ w44734;
	assign w32520 = w32615 ^ w32564;
	assign w32602 = w47835 ^ w32520;
	assign w32600 = w32601 & w32602;
	assign w32598 = w32606 ^ w32600;
	assign w32519 = w32600 ^ w32564;
	assign w32518 = w32600 ^ w32617;
	assign w32513 = w32518 ^ w32614;
	assign w32524 = w32550 ^ w44734;
	assign w32608 = w32524 ^ w32549;
	assign w32599 = w32600 ^ w32608;
	assign w32605 = w32606 ^ w32608;
	assign w32604 = w32607 & w32605;
	assign w32603 = w32604 ^ w32566;
	assign w32515 = w32604 ^ w32616;
	assign w32511 = w32515 ^ w32551;
	assign w32514 = w47829 ^ w32511;
	assign w32591 = w32513 ^ w32514;
	assign w32512 = w32604 ^ w32560;
	assign w32510 = w47831 ^ w32511;
	assign w32597 = w32608 & w32598;
	assign w32595 = w32597 ^ w32605;
	assign w32594 = w32603 & w32595;
	assign w32559 = w32594 ^ w32569;
	assign w32593 = w32559 ^ w32561;
	assign w32517 = w32594 ^ w32618;
	assign w32590 = w32559 ^ w32512;
	assign w32585 = w32599 & w47836;
	assign w32584 = w32590 & w32620;
	assign w32583 = w32593 & w32632;
	assign w32582 = w32603 & w32622;
	assign w32526 = w32582 ^ w32583;
	assign w32581 = w32591 & w32623;
	assign w32576 = w32599 & w32631;
	assign w32575 = w32590 & w32635;
	assign w32542 = w32584 ^ w32575;
	assign w32574 = w32593 & w32628;
	assign w32544 = w32582 ^ w32574;
	assign w32573 = w32603 & w32629;
	assign w32572 = w32591 & w32634;
	assign w44735 = w32583 ^ w32584;
	assign w44737 = w32597 ^ w32615;
	assign w32556 = w47835 ^ w44737;
	assign w32596 = w32556 ^ w32519;
	assign w32509 = w32556 ^ w32517;
	assign w32516 = w32546 ^ w32509;
	assign w32592 = w32513 ^ w32516;
	assign w32588 = w32509 ^ w32510;
	assign w32586 = w32596 & w32625;
	assign w32580 = w32588 & w32621;
	assign w32541 = w32580 ^ w32583;
	assign w32538 = ~w32541;
	assign w32537 = w32580 ^ w32581;
	assign w32579 = w32592 & w32624;
	assign w32577 = w32596 & w32627;
	assign w32557 = w32575 ^ w32579;
	assign w32535 = ~w32557;
	assign w32534 = w32535 ^ w32573;
	assign w32571 = w32588 & w32636;
	assign w32570 = w32592 & w32633;
	assign w32536 = w32581 ^ w32570;
	assign w32532 = ~w32536;
	assign w43590 = w32571 ^ w32572;
	assign w32540 = w32544 ^ w43590;
	assign w32539 = w32535 ^ w32540;
	assign w32639 = w32538 ^ w32539;
	assign w32553 = w32577 ^ w43590;
	assign w32565 = w32580 ^ w44735;
	assign w32531 = w32576 ^ w32565;
	assign w32528 = ~w32531;
	assign w32525 = w32581 ^ w32565;
	assign w32589 = w44737 ^ w32567;
	assign w32587 = w32589 & w32626;
	assign w32578 = w32589 & w32630;
	assign w32554 = w32578 ^ w32553;
	assign w32558 = w32586 ^ w32554;
	assign w32563 = w32587 ^ w32558;
	assign w48472 = w44735 ^ w32563;
	assign w6010 = w48468 ^ w48472;
	assign w6136 = w6134 ^ w6010;
	assign w6260 = w6258 ^ w48472;
	assign w5949 = w6260 ^ w6259;
	assign w48361 = w5949 ^ w6002;
	assign w47712 = w48361 ^ w52;
	assign w32638 = w32563 ^ w32537;
	assign w32527 = w32585 ^ w32558;
	assign w48471 = w32526 ^ w32527;
	assign w6005 = w48467 ^ w48471;
	assign w6133 = w6142 ^ w6005;
	assign w6163 = w6160 ^ w6005;
	assign w6262 = w6023 ^ w48471;
	assign w5948 = w6262 ^ w6261;
	assign w48360 = w5948 ^ w5998;
	assign w47713 = w48360 ^ w51;
	assign w48473 = w32554 ^ w32525;
	assign w6031 = w48469 ^ w48473;
	assign w6021 = w48460 ^ w48473;
	assign w6155 = w6031 ^ w48467;
	assign w6162 = w6031 ^ w6161;
	assign w48369 = w6163 ^ w6162;
	assign w47704 = w48369 ^ w60;
	assign w6270 = w6021 ^ w48471;
	assign w5944 = w6270 ^ w6269;
	assign w48345 = w5944 ^ w6010;
	assign w47728 = w48345 ^ w36;
	assign w6274 = ~w6021;
	assign w44736 = w32585 ^ w32587;
	assign w32543 = w44736 ^ w32540;
	assign w32640 = w32542 ^ w32543;
	assign w32530 = w32534 ^ w44736;
	assign w32533 = w32572 ^ w32530;
	assign w32637 = w32532 ^ w32533;
	assign w32529 = w32553 ^ w32530;
	assign w48470 = w32528 ^ w32529;
	assign w6000 = w48466 ^ w48470;
	assign w6144 = w6142 ^ w48470;
	assign w6156 = w5998 ^ w6000;
	assign w48368 = w6156 ^ w6155;
	assign w47705 = w48368 ^ w59;
	assign w6273 = w6274 ^ w48470;
	assign w5943 = w6273 ^ w6272;
	assign w48344 = w5943 ^ w6005;
	assign w47729 = w48344 ^ w35;
	assign w44857 = w35559 ^ w35562;
	assign w35472 = w35498 ^ w44857;
	assign w35556 = w35472 ^ w35497;
	assign w35553 = w35554 ^ w35556;
	assign w35512 = w35560 ^ w44857;
	assign w35468 = w35563 ^ w35512;
	assign w35550 = w1701 ^ w35468;
	assign w44860 = w35559 ^ w35565;
	assign w35471 = w35503 ^ w44860;
	assign w35514 = w1705 ^ w35471;
	assign w35549 = w35554 ^ w35514;
	assign w35548 = w35549 & w35550;
	assign w35547 = w35548 ^ w35556;
	assign w35546 = w35554 ^ w35548;
	assign w35467 = w35548 ^ w35512;
	assign w35466 = w35548 ^ w35565;
	assign w35461 = w35466 ^ w35562;
	assign w35545 = w35556 & w35546;
	assign w35543 = w35545 ^ w35553;
	assign w35533 = w35547 & w1700;
	assign w35524 = w35547 & w35579;
	assign w44859 = w35545 ^ w35563;
	assign w35537 = w44859 ^ w35515;
	assign w35535 = w35537 & w35574;
	assign w35526 = w35537 & w35578;
	assign w35504 = w1701 ^ w44859;
	assign w35544 = w35504 ^ w35467;
	assign w35534 = w35544 & w35573;
	assign w35525 = w35544 & w35575;
	assign w35509 = w44860 ^ w35494;
	assign w35555 = w35517 ^ w35509;
	assign w35552 = w35555 & w35553;
	assign w35551 = w35552 ^ w35514;
	assign w35463 = w35552 ^ w35564;
	assign w35459 = w35463 ^ w35499;
	assign w35462 = w1707 ^ w35459;
	assign w35539 = w35461 ^ w35462;
	assign w35460 = w35552 ^ w35508;
	assign w35458 = w1705 ^ w35459;
	assign w35542 = w35551 & w35543;
	assign w35507 = w35542 ^ w35517;
	assign w35541 = w35507 ^ w35509;
	assign w35465 = w35542 ^ w35566;
	assign w35457 = w35504 ^ w35465;
	assign w35464 = w35494 ^ w35457;
	assign w35540 = w35461 ^ w35464;
	assign w35538 = w35507 ^ w35460;
	assign w35536 = w35457 ^ w35458;
	assign w35532 = w35538 & w35568;
	assign w35531 = w35541 & w35580;
	assign w35530 = w35551 & w35570;
	assign w35474 = w35530 ^ w35531;
	assign w35529 = w35539 & w35571;
	assign w35528 = w35536 & w35569;
	assign w35489 = w35528 ^ w35531;
	assign w35486 = ~w35489;
	assign w35485 = w35528 ^ w35529;
	assign w35527 = w35540 & w35572;
	assign w35523 = w35538 & w35583;
	assign w35505 = w35523 ^ w35527;
	assign w35490 = w35532 ^ w35523;
	assign w35483 = ~w35505;
	assign w35522 = w35541 & w35576;
	assign w35492 = w35530 ^ w35522;
	assign w35521 = w35551 & w35577;
	assign w35482 = w35483 ^ w35521;
	assign w35520 = w35539 & w35582;
	assign w35519 = w35536 & w35584;
	assign w35518 = w35540 & w35581;
	assign w35484 = w35529 ^ w35518;
	assign w35480 = ~w35484;
	assign w44858 = w35519 ^ w35520;
	assign w35501 = w35525 ^ w44858;
	assign w35502 = w35526 ^ w35501;
	assign w35506 = w35534 ^ w35502;
	assign w35511 = w35535 ^ w35506;
	assign w35586 = w35511 ^ w35485;
	assign w35475 = w35533 ^ w35506;
	assign w48040 = w35474 ^ w35475;
	assign w48043 = ~w35586;
	assign w35488 = w35492 ^ w44858;
	assign w35487 = w35483 ^ w35488;
	assign w35587 = w35486 ^ w35487;
	assign w48038 = ~w35587;
	assign w44861 = w35531 ^ w35532;
	assign w48041 = w44861 ^ w35511;
	assign w35513 = w35528 ^ w44861;
	assign w35479 = w35524 ^ w35513;
	assign w35476 = ~w35479;
	assign w35473 = w35529 ^ w35513;
	assign w48044 = w35502 ^ w35473;
	assign w44862 = w35533 ^ w35535;
	assign w35491 = w44862 ^ w35488;
	assign w35588 = w35490 ^ w35491;
	assign w48037 = ~w35588;
	assign w35478 = w35482 ^ w44862;
	assign w35481 = w35520 ^ w35478;
	assign w35585 = w35480 ^ w35481;
	assign w35477 = w35501 ^ w35478;
	assign w48039 = w35476 ^ w35477;
	assign w48042 = ~w35585;
	assign w44868 = w35827 ^ w35833;
	assign w35739 = w35771 ^ w44868;
	assign w35782 = w1450 ^ w35739;
	assign w35817 = w35822 ^ w35782;
	assign w35777 = w44868 ^ w35762;
	assign w35823 = w35785 ^ w35777;
	assign w44869 = w35827 ^ w35830;
	assign w35780 = w35828 ^ w44869;
	assign w35736 = w35831 ^ w35780;
	assign w35818 = w1446 ^ w35736;
	assign w35816 = w35817 & w35818;
	assign w35814 = w35822 ^ w35816;
	assign w35734 = w35816 ^ w35833;
	assign w35729 = w35734 ^ w35830;
	assign w35735 = w35816 ^ w35780;
	assign w35740 = w35766 ^ w44869;
	assign w35824 = w35740 ^ w35765;
	assign w35815 = w35816 ^ w35824;
	assign w35821 = w35822 ^ w35824;
	assign w35820 = w35823 & w35821;
	assign w35819 = w35820 ^ w35782;
	assign w35731 = w35820 ^ w35832;
	assign w35727 = w35731 ^ w35767;
	assign w35730 = w1452 ^ w35727;
	assign w35807 = w35729 ^ w35730;
	assign w35728 = w35820 ^ w35776;
	assign w35726 = w1450 ^ w35727;
	assign w35813 = w35824 & w35814;
	assign w35811 = w35813 ^ w35821;
	assign w35810 = w35819 & w35811;
	assign w35775 = w35810 ^ w35785;
	assign w35809 = w35775 ^ w35777;
	assign w35733 = w35810 ^ w35834;
	assign w35806 = w35775 ^ w35728;
	assign w35801 = w35815 & w1445;
	assign w35800 = w35806 & w35836;
	assign w35799 = w35809 & w35848;
	assign w35798 = w35819 & w35838;
	assign w35742 = w35798 ^ w35799;
	assign w35797 = w35807 & w35839;
	assign w35792 = w35815 & w35847;
	assign w35791 = w35806 & w35851;
	assign w35758 = w35800 ^ w35791;
	assign w35790 = w35809 & w35844;
	assign w35760 = w35798 ^ w35790;
	assign w35789 = w35819 & w35845;
	assign w35788 = w35807 & w35850;
	assign w44871 = w35799 ^ w35800;
	assign w44873 = w35813 ^ w35831;
	assign w35805 = w44873 ^ w35783;
	assign w35794 = w35805 & w35846;
	assign w35803 = w35805 & w35842;
	assign w44872 = w35801 ^ w35803;
	assign w35772 = w1446 ^ w44873;
	assign w35812 = w35772 ^ w35735;
	assign w35725 = w35772 ^ w35733;
	assign w35732 = w35762 ^ w35725;
	assign w35808 = w35729 ^ w35732;
	assign w35804 = w35725 ^ w35726;
	assign w35802 = w35812 & w35841;
	assign w35796 = w35804 & w35837;
	assign w35781 = w35796 ^ w44871;
	assign w35757 = w35796 ^ w35799;
	assign w35754 = ~w35757;
	assign w35753 = w35796 ^ w35797;
	assign w35747 = w35792 ^ w35781;
	assign w35744 = ~w35747;
	assign w35741 = w35797 ^ w35781;
	assign w35795 = w35808 & w35840;
	assign w35773 = w35791 ^ w35795;
	assign w35751 = ~w35773;
	assign w35750 = w35751 ^ w35789;
	assign w35746 = w35750 ^ w44872;
	assign w35749 = w35788 ^ w35746;
	assign w35793 = w35812 & w35843;
	assign w35787 = w35804 & w35852;
	assign w35786 = w35808 & w35849;
	assign w35752 = w35797 ^ w35786;
	assign w35748 = ~w35752;
	assign w35853 = w35748 ^ w35749;
	assign w47978 = ~w35853;
	assign w1490 = w1904 ^ w47978;
	assign w1521 = w1935 ^ w1490;
	assign w1553 = w1967 ^ w1521;
	assign w1585 = w1999 ^ w1553;
	assign w1745 = w1490 ^ w48042;
	assign w1776 = w1521 ^ w1745;
	assign w1808 = w1553 ^ w1776;
	assign w1840 = w1585 ^ w1808;
	assign w44870 = w35787 ^ w35788;
	assign w35769 = w35793 ^ w44870;
	assign w35745 = w35769 ^ w35746;
	assign w47975 = w35744 ^ w35745;
	assign w1487 = w1901 ^ w47975;
	assign w1518 = w1932 ^ w1487;
	assign w1550 = w1964 ^ w1518;
	assign w1582 = w1996 ^ w1550;
	assign w1742 = w1487 ^ w48039;
	assign w1773 = w1518 ^ w1742;
	assign w1805 = w1550 ^ w1773;
	assign w1837 = w1582 ^ w1805;
	assign w35770 = w35794 ^ w35769;
	assign w47980 = w35770 ^ w35741;
	assign w1492 = w1906 ^ w47980;
	assign w1523 = w1937 ^ w1492;
	assign w1555 = w1969 ^ w1523;
	assign w1587 = w2001 ^ w1555;
	assign w1747 = w1492 ^ w48044;
	assign w1778 = w1523 ^ w1747;
	assign w1810 = w1555 ^ w1778;
	assign w1842 = w1587 ^ w1810;
	assign w35447 = w1842 ^ w1837;
	assign w35715 = w1587 ^ w1582;
	assign w35360 = w1840 ^ w1842;
	assign w35628 = w1585 ^ w1587;
	assign w35774 = w35802 ^ w35770;
	assign w35779 = w35803 ^ w35774;
	assign w35854 = w35779 ^ w35753;
	assign w47979 = ~w35854;
	assign w1491 = w1905 ^ w47979;
	assign w1522 = w1936 ^ w1491;
	assign w1554 = w1968 ^ w1522;
	assign w1586 = w2000 ^ w1554;
	assign w1746 = w1491 ^ w48043;
	assign w1777 = w1522 ^ w1746;
	assign w1809 = w1554 ^ w1777;
	assign w1841 = w1586 ^ w1809;
	assign w47977 = w44871 ^ w35779;
	assign w1489 = w1903 ^ w47977;
	assign w1744 = w1489 ^ w48041;
	assign w1520 = w1934 ^ w1489;
	assign w1775 = w1520 ^ w1744;
	assign w1552 = w1966 ^ w1520;
	assign w1584 = w1998 ^ w1552;
	assign w35716 = w1584 ^ w1587;
	assign w35718 = w1582 ^ w1584;
	assign w1807 = w1552 ^ w1775;
	assign w35630 = w1584 ^ w1586;
	assign w1839 = w1584 ^ w1807;
	assign w35448 = w1839 ^ w1842;
	assign w35362 = w1839 ^ w1841;
	assign w35450 = w1837 ^ w1839;
	assign w35743 = w35801 ^ w35774;
	assign w35435 = w35360 ^ w35450;
	assign w35322 = w35362 ^ w35360;
	assign w35321 = w35362 ^ w1840;
	assign w35426 = w35450 & w35435;
	assign w47976 = w35742 ^ w35743;
	assign w35703 = w35628 ^ w35718;
	assign w35590 = w35630 ^ w35628;
	assign w35589 = w35630 ^ w1585;
	assign w35694 = w35718 & w35703;
	assign w1488 = w1902 ^ w47976;
	assign w1519 = w1933 ^ w1488;
	assign w1743 = w1488 ^ w48040;
	assign w1774 = w1519 ^ w1743;
	assign w1551 = w1965 ^ w1519;
	assign w1583 = w1997 ^ w1551;
	assign w1806 = w1551 ^ w1774;
	assign w1838 = w1583 ^ w1806;
	assign w35336 = w1838 ^ w1837;
	assign w35604 = w1583 ^ w1582;
	assign w35756 = w35760 ^ w44870;
	assign w35759 = w44872 ^ w35756;
	assign w35856 = w35758 ^ w35759;
	assign w35755 = w35751 ^ w35756;
	assign w35855 = w35754 ^ w35755;
	assign w47973 = ~w35856;
	assign w1485 = w1899 ^ w47973;
	assign w1516 = w1930 ^ w1485;
	assign w1548 = w1962 ^ w1516;
	assign w1580 = w1994 ^ w1548;
	assign w1740 = w1485 ^ w48037;
	assign w1771 = w1516 ^ w1740;
	assign w1803 = w1548 ^ w1771;
	assign w1835 = w1580 ^ w1803;
	assign w35366 = w1835 ^ w1841;
	assign w35443 = w35360 ^ w35366;
	assign w35446 = w1840 ^ w35366;
	assign w35445 = w1835 ^ w35321;
	assign w35431 = w35445 & w1835;
	assign w35634 = w1580 ^ w1586;
	assign w35711 = w35628 ^ w35634;
	assign w35714 = w1585 ^ w35634;
	assign w35713 = w1580 ^ w35589;
	assign w35699 = w35713 & w1580;
	assign w47974 = ~w35855;
	assign w1486 = w1900 ^ w47974;
	assign w1517 = w1931 ^ w1486;
	assign w1549 = w1963 ^ w1517;
	assign w1581 = w1995 ^ w1549;
	assign w1741 = w1486 ^ w48038;
	assign w1772 = w1517 ^ w1741;
	assign w1804 = w1549 ^ w1772;
	assign w1836 = w1581 ^ w1804;
	assign w35359 = w1836 ^ w1838;
	assign w35361 = w1837 ^ w35359;
	assign w35437 = w1841 ^ w35361;
	assign w35434 = w1840 ^ w35361;
	assign w35436 = w35366 ^ w35361;
	assign w35442 = w1836 ^ w35446;
	assign w35440 = w35359 ^ w35448;
	assign w35439 = w1835 ^ w35440;
	assign w35376 = w1836 ^ w1837;
	assign w35441 = w35376 ^ w35443;
	assign w35444 = w35448 ^ w35376;
	assign w35438 = w35359 ^ w35322;
	assign w35449 = w1842 ^ w1836;
	assign w35433 = w35440 & w35444;
	assign w35365 = w35433 ^ w35362;
	assign w35432 = w35441 & w35439;
	assign w35383 = w35426 ^ w35432;
	assign w35430 = w35449 & w35434;
	assign w35364 = w35430 ^ w35360;
	assign w35429 = w35446 & w35442;
	assign w35428 = w35443 & w35436;
	assign w35427 = w35448 & w35437;
	assign w35363 = w35427 ^ w35361;
	assign w35369 = w35365 ^ w35363;
	assign w35374 = w1842 ^ w35369;
	assign w35424 = w35383 ^ w35374;
	assign w35335 = w35426 ^ w35427;
	assign w35382 = w35335 ^ w35336;
	assign w35381 = w35382 ^ w35364;
	assign w35423 = w35429 ^ w35381;
	assign w35425 = w35447 & w35438;
	assign w35420 = w35424 & w35423;
	assign w35627 = w1581 ^ w1583;
	assign w35629 = w1582 ^ w35627;
	assign w35705 = w1586 ^ w35629;
	assign w35702 = w1585 ^ w35629;
	assign w35704 = w35634 ^ w35629;
	assign w35710 = w1581 ^ w35714;
	assign w35708 = w35627 ^ w35716;
	assign w35707 = w1580 ^ w35708;
	assign w35644 = w1581 ^ w1582;
	assign w35709 = w35644 ^ w35711;
	assign w35712 = w35716 ^ w35644;
	assign w35706 = w35627 ^ w35590;
	assign w35717 = w1587 ^ w1581;
	assign w35701 = w35708 & w35712;
	assign w35633 = w35701 ^ w35630;
	assign w35700 = w35709 & w35707;
	assign w35651 = w35694 ^ w35700;
	assign w35698 = w35717 & w35702;
	assign w35632 = w35698 ^ w35628;
	assign w35697 = w35714 & w35710;
	assign w35696 = w35711 & w35704;
	assign w35695 = w35716 & w35705;
	assign w35631 = w35695 ^ w35629;
	assign w35637 = w35633 ^ w35631;
	assign w35642 = w1587 ^ w35637;
	assign w35692 = w35651 ^ w35642;
	assign w35603 = w35694 ^ w35695;
	assign w35650 = w35603 ^ w35604;
	assign w35649 = w35650 ^ w35632;
	assign w35691 = w35697 ^ w35649;
	assign w35693 = w35715 & w35706;
	assign w35688 = w35692 & w35691;
	assign w44851 = w35425 ^ w35431;
	assign w35337 = w35369 ^ w44851;
	assign w35380 = w1840 ^ w35337;
	assign w35415 = w35420 ^ w35380;
	assign w35375 = w44851 ^ w35360;
	assign w35421 = w35383 ^ w35375;
	assign w44852 = w35425 ^ w35428;
	assign w35378 = w35426 ^ w44852;
	assign w35334 = w35429 ^ w35378;
	assign w35416 = w1836 ^ w35334;
	assign w35414 = w35415 & w35416;
	assign w35412 = w35420 ^ w35414;
	assign w35333 = w35414 ^ w35378;
	assign w35332 = w35414 ^ w35431;
	assign w35327 = w35332 ^ w35428;
	assign w35338 = w35364 ^ w44852;
	assign w35422 = w35338 ^ w35363;
	assign w35413 = w35414 ^ w35422;
	assign w35419 = w35420 ^ w35422;
	assign w35418 = w35421 & w35419;
	assign w35417 = w35418 ^ w35380;
	assign w35329 = w35418 ^ w35430;
	assign w35325 = w35329 ^ w35365;
	assign w35328 = w1842 ^ w35325;
	assign w35405 = w35327 ^ w35328;
	assign w35326 = w35418 ^ w35374;
	assign w35324 = w1840 ^ w35325;
	assign w35411 = w35422 & w35412;
	assign w35409 = w35411 ^ w35419;
	assign w35408 = w35417 & w35409;
	assign w35373 = w35408 ^ w35383;
	assign w35407 = w35373 ^ w35375;
	assign w35331 = w35408 ^ w35432;
	assign w35404 = w35373 ^ w35326;
	assign w35399 = w35413 & w1835;
	assign w35398 = w35404 & w35434;
	assign w35397 = w35407 & w35446;
	assign w35396 = w35417 & w35436;
	assign w35340 = w35396 ^ w35397;
	assign w35395 = w35405 & w35437;
	assign w35390 = w35413 & w35445;
	assign w35389 = w35404 & w35449;
	assign w35356 = w35398 ^ w35389;
	assign w35388 = w35407 & w35442;
	assign w35358 = w35396 ^ w35388;
	assign w35387 = w35417 & w35443;
	assign w35386 = w35405 & w35448;
	assign w44854 = w35397 ^ w35398;
	assign w44856 = w35411 ^ w35429;
	assign w35403 = w44856 ^ w35381;
	assign w35401 = w35403 & w35440;
	assign w35392 = w35403 & w35444;
	assign w44855 = w35399 ^ w35401;
	assign w35370 = w1836 ^ w44856;
	assign w35410 = w35370 ^ w35333;
	assign w35323 = w35370 ^ w35331;
	assign w35330 = w35360 ^ w35323;
	assign w35406 = w35327 ^ w35330;
	assign w35402 = w35323 ^ w35324;
	assign w35400 = w35410 & w35439;
	assign w35394 = w35402 & w35435;
	assign w35379 = w35394 ^ w44854;
	assign w35355 = w35394 ^ w35397;
	assign w35352 = ~w35355;
	assign w35351 = w35394 ^ w35395;
	assign w35345 = w35390 ^ w35379;
	assign w35342 = ~w35345;
	assign w35339 = w35395 ^ w35379;
	assign w35393 = w35406 & w35438;
	assign w35371 = w35389 ^ w35393;
	assign w35349 = ~w35371;
	assign w35348 = w35349 ^ w35387;
	assign w35344 = w35348 ^ w44855;
	assign w35347 = w35386 ^ w35344;
	assign w35391 = w35410 & w35441;
	assign w35385 = w35402 & w35450;
	assign w35384 = w35406 & w35447;
	assign w35350 = w35395 ^ w35384;
	assign w35346 = ~w35350;
	assign w35451 = w35346 ^ w35347;
	assign w48074 = ~w35451;
	assign w44853 = w35385 ^ w35386;
	assign w35367 = w35391 ^ w44853;
	assign w35368 = w35392 ^ w35367;
	assign w35372 = w35400 ^ w35368;
	assign w35377 = w35401 ^ w35372;
	assign w48073 = w44854 ^ w35377;
	assign w35452 = w35377 ^ w35351;
	assign w35343 = w35367 ^ w35344;
	assign w48071 = w35342 ^ w35343;
	assign w35341 = w35399 ^ w35372;
	assign w48072 = w35340 ^ w35341;
	assign w48076 = w35368 ^ w35339;
	assign w48075 = ~w35452;
	assign w35354 = w35358 ^ w44853;
	assign w35357 = w44855 ^ w35354;
	assign w35454 = w35356 ^ w35357;
	assign w35353 = w35349 ^ w35354;
	assign w35453 = w35352 ^ w35353;
	assign w48069 = ~w35454;
	assign w48070 = ~w35453;
	assign w44863 = w35693 ^ w35699;
	assign w35643 = w44863 ^ w35628;
	assign w35689 = w35651 ^ w35643;
	assign w35605 = w35637 ^ w44863;
	assign w35648 = w1585 ^ w35605;
	assign w35683 = w35688 ^ w35648;
	assign w44864 = w35693 ^ w35696;
	assign w35646 = w35694 ^ w44864;
	assign w35602 = w35697 ^ w35646;
	assign w35684 = w1581 ^ w35602;
	assign w35682 = w35683 & w35684;
	assign w35680 = w35688 ^ w35682;
	assign w35601 = w35682 ^ w35646;
	assign w35600 = w35682 ^ w35699;
	assign w35595 = w35600 ^ w35696;
	assign w35606 = w35632 ^ w44864;
	assign w35690 = w35606 ^ w35631;
	assign w35681 = w35682 ^ w35690;
	assign w35687 = w35688 ^ w35690;
	assign w35686 = w35689 & w35687;
	assign w35685 = w35686 ^ w35648;
	assign w35597 = w35686 ^ w35698;
	assign w35593 = w35597 ^ w35633;
	assign w35596 = w1587 ^ w35593;
	assign w35673 = w35595 ^ w35596;
	assign w35594 = w35686 ^ w35642;
	assign w35592 = w1585 ^ w35593;
	assign w35679 = w35690 & w35680;
	assign w35677 = w35679 ^ w35687;
	assign w35676 = w35685 & w35677;
	assign w35641 = w35676 ^ w35651;
	assign w35675 = w35641 ^ w35643;
	assign w35599 = w35676 ^ w35700;
	assign w35672 = w35641 ^ w35594;
	assign w35667 = w35681 & w1580;
	assign w35666 = w35672 & w35702;
	assign w35665 = w35675 & w35714;
	assign w35664 = w35685 & w35704;
	assign w35608 = w35664 ^ w35665;
	assign w35663 = w35673 & w35705;
	assign w35658 = w35681 & w35713;
	assign w35657 = w35672 & w35717;
	assign w35624 = w35666 ^ w35657;
	assign w35656 = w35675 & w35710;
	assign w35626 = w35664 ^ w35656;
	assign w35655 = w35685 & w35711;
	assign w35654 = w35673 & w35716;
	assign w44865 = w35665 ^ w35666;
	assign w44867 = w35679 ^ w35697;
	assign w35638 = w1581 ^ w44867;
	assign w35678 = w35638 ^ w35601;
	assign w35668 = w35678 & w35707;
	assign w35659 = w35678 & w35709;
	assign w35591 = w35638 ^ w35599;
	assign w35670 = w35591 ^ w35592;
	assign w35662 = w35670 & w35703;
	assign w35623 = w35662 ^ w35665;
	assign w35620 = ~w35623;
	assign w35619 = w35662 ^ w35663;
	assign w35653 = w35670 & w35718;
	assign w43598 = w35653 ^ w35654;
	assign w35622 = w35626 ^ w43598;
	assign w35635 = w35659 ^ w43598;
	assign w35598 = w35628 ^ w35591;
	assign w35647 = w35662 ^ w44865;
	assign w35613 = w35658 ^ w35647;
	assign w35610 = ~w35613;
	assign w35607 = w35663 ^ w35647;
	assign w35674 = w35595 ^ w35598;
	assign w35652 = w35674 & w35715;
	assign w35618 = w35663 ^ w35652;
	assign w35614 = ~w35618;
	assign w35661 = w35674 & w35706;
	assign w35639 = w35657 ^ w35661;
	assign w35617 = ~w35639;
	assign w35621 = w35617 ^ w35622;
	assign w35721 = w35620 ^ w35621;
	assign w48006 = ~w35721;
	assign w1613 = w2027 ^ w48006;
	assign w1645 = w1390 ^ w1613;
	assign w1677 = w1422 ^ w1645;
	assign w1709 = w1454 ^ w1677;
	assign w1868 = w1613 ^ w48070;
	assign w880 = w1645 ^ w1868;
	assign w912 = w1677 ^ w880;
	assign w944 = w1709 ^ w912;
	assign w35616 = w35617 ^ w35655;
	assign w35671 = w44867 ^ w35649;
	assign w35669 = w35671 & w35708;
	assign w35660 = w35671 & w35712;
	assign w35636 = w35660 ^ w35635;
	assign w35640 = w35668 ^ w35636;
	assign w35645 = w35669 ^ w35640;
	assign w48009 = w44865 ^ w35645;
	assign w1616 = w2030 ^ w48009;
	assign w1648 = w1393 ^ w1616;
	assign w1680 = w1425 ^ w1648;
	assign w1712 = w1457 ^ w1680;
	assign w1871 = w1616 ^ w48073;
	assign w883 = w1648 ^ w1871;
	assign w915 = w1680 ^ w883;
	assign w947 = w1712 ^ w915;
	assign w35720 = w35645 ^ w35619;
	assign w35609 = w35667 ^ w35640;
	assign w48008 = w35608 ^ w35609;
	assign w1615 = w2029 ^ w48008;
	assign w1647 = w1392 ^ w1615;
	assign w1679 = w1424 ^ w1647;
	assign w1711 = w1456 ^ w1679;
	assign w1870 = w1615 ^ w48072;
	assign w882 = w1647 ^ w1870;
	assign w914 = w1679 ^ w882;
	assign w946 = w1711 ^ w914;
	assign w48012 = w35636 ^ w35607;
	assign w1619 = w2033 ^ w48012;
	assign w1651 = w1396 ^ w1619;
	assign w1683 = w1428 ^ w1651;
	assign w1715 = w1460 ^ w1683;
	assign w1874 = w1619 ^ w48076;
	assign w886 = w1651 ^ w1874;
	assign w918 = w1683 ^ w886;
	assign w950 = w1715 ^ w918;
	assign w48011 = ~w35720;
	assign w1618 = w2032 ^ w48011;
	assign w1650 = w1395 ^ w1618;
	assign w1682 = w1427 ^ w1650;
	assign w1714 = w1459 ^ w1682;
	assign w1873 = w1618 ^ w48075;
	assign w885 = w1650 ^ w1873;
	assign w917 = w1682 ^ w885;
	assign w949 = w1714 ^ w917;
	assign w38039 = w944 ^ w946;
	assign w38042 = w947 ^ w949;
	assign w38128 = w947 ^ w950;
	assign w38120 = w38039 ^ w38128;
	assign w38129 = w950 ^ w944;
	assign w38307 = w1709 ^ w1711;
	assign w38310 = w1712 ^ w1714;
	assign w38396 = w1712 ^ w1715;
	assign w38388 = w38307 ^ w38396;
	assign w38397 = w1715 ^ w1709;
	assign w44866 = w35667 ^ w35669;
	assign w35625 = w44866 ^ w35622;
	assign w35722 = w35624 ^ w35625;
	assign w48005 = ~w35722;
	assign w1612 = w2026 ^ w48005;
	assign w1644 = w1389 ^ w1612;
	assign w1676 = w1421 ^ w1644;
	assign w1708 = w1453 ^ w1676;
	assign w38314 = w1708 ^ w1714;
	assign w38387 = w1708 ^ w38388;
	assign w1867 = w1612 ^ w48069;
	assign w879 = w1644 ^ w1867;
	assign w911 = w1676 ^ w879;
	assign w943 = w1708 ^ w911;
	assign w38046 = w943 ^ w949;
	assign w38119 = w943 ^ w38120;
	assign w35612 = w35616 ^ w44866;
	assign w35615 = w35654 ^ w35612;
	assign w35719 = w35614 ^ w35615;
	assign w35611 = w35635 ^ w35612;
	assign w48007 = w35610 ^ w35611;
	assign w1614 = w2028 ^ w48007;
	assign w1646 = w1391 ^ w1614;
	assign w1678 = w1423 ^ w1646;
	assign w1710 = w1455 ^ w1678;
	assign w1869 = w1614 ^ w48071;
	assign w881 = w1646 ^ w1869;
	assign w913 = w1678 ^ w881;
	assign w945 = w1710 ^ w913;
	assign w48010 = ~w35719;
	assign w1617 = w2031 ^ w48010;
	assign w1649 = w1394 ^ w1617;
	assign w1681 = w1426 ^ w1649;
	assign w1713 = w1458 ^ w1681;
	assign w1872 = w1617 ^ w48074;
	assign w884 = w1649 ^ w1872;
	assign w916 = w1681 ^ w884;
	assign w948 = w1713 ^ w916;
	assign w38040 = w948 ^ w950;
	assign w38041 = w945 ^ w38039;
	assign w38117 = w949 ^ w38041;
	assign w38114 = w948 ^ w38041;
	assign w38116 = w38046 ^ w38041;
	assign w38123 = w38040 ^ w38046;
	assign w38056 = w944 ^ w945;
	assign w38121 = w38056 ^ w38123;
	assign w38124 = w38128 ^ w38056;
	assign w38130 = w945 ^ w947;
	assign w38115 = w38040 ^ w38130;
	assign w38126 = w948 ^ w38046;
	assign w38122 = w944 ^ w38126;
	assign w38016 = w946 ^ w945;
	assign w38002 = w38042 ^ w38040;
	assign w38118 = w38039 ^ w38002;
	assign w38001 = w38042 ^ w948;
	assign w38125 = w943 ^ w38001;
	assign w38127 = w950 ^ w945;
	assign w38113 = w38120 & w38124;
	assign w38045 = w38113 ^ w38042;
	assign w38112 = w38121 & w38119;
	assign w38111 = w38125 & w943;
	assign w38110 = w38129 & w38114;
	assign w38044 = w38110 ^ w38040;
	assign w38109 = w38126 & w38122;
	assign w38108 = w38123 & w38116;
	assign w38107 = w38128 & w38117;
	assign w38043 = w38107 ^ w38041;
	assign w38049 = w38045 ^ w38043;
	assign w38054 = w950 ^ w38049;
	assign w38106 = w38130 & w38115;
	assign w38063 = w38106 ^ w38112;
	assign w38104 = w38063 ^ w38054;
	assign w38015 = w38106 ^ w38107;
	assign w38062 = w38015 ^ w38016;
	assign w38061 = w38062 ^ w38044;
	assign w38103 = w38109 ^ w38061;
	assign w38105 = w38127 & w38118;
	assign w38100 = w38104 & w38103;
	assign w38308 = w1713 ^ w1715;
	assign w38309 = w1710 ^ w38307;
	assign w38385 = w1714 ^ w38309;
	assign w38382 = w1713 ^ w38309;
	assign w38384 = w38314 ^ w38309;
	assign w38391 = w38308 ^ w38314;
	assign w38324 = w1709 ^ w1710;
	assign w38389 = w38324 ^ w38391;
	assign w38392 = w38396 ^ w38324;
	assign w38398 = w1710 ^ w1712;
	assign w38383 = w38308 ^ w38398;
	assign w38394 = w1713 ^ w38314;
	assign w38390 = w1709 ^ w38394;
	assign w38284 = w1711 ^ w1710;
	assign w38270 = w38310 ^ w38308;
	assign w38386 = w38307 ^ w38270;
	assign w38269 = w38310 ^ w1713;
	assign w38393 = w1708 ^ w38269;
	assign w38395 = w1715 ^ w1710;
	assign w38381 = w38388 & w38392;
	assign w38313 = w38381 ^ w38310;
	assign w38380 = w38389 & w38387;
	assign w38379 = w38393 & w1708;
	assign w38378 = w38397 & w38382;
	assign w38312 = w38378 ^ w38308;
	assign w38377 = w38394 & w38390;
	assign w38376 = w38391 & w38384;
	assign w38375 = w38396 & w38385;
	assign w38311 = w38375 ^ w38309;
	assign w38317 = w38313 ^ w38311;
	assign w38322 = w1715 ^ w38317;
	assign w38374 = w38398 & w38383;
	assign w38331 = w38374 ^ w38380;
	assign w38372 = w38331 ^ w38322;
	assign w38283 = w38374 ^ w38375;
	assign w38330 = w38283 ^ w38284;
	assign w38329 = w38330 ^ w38312;
	assign w38371 = w38377 ^ w38329;
	assign w38373 = w38395 & w38386;
	assign w38368 = w38372 & w38371;
	assign w44880 = w36095 ^ w36101;
	assign w36045 = w44880 ^ w36030;
	assign w36091 = w36053 ^ w36045;
	assign w36007 = w36039 ^ w44880;
	assign w36050 = w47815 ^ w36007;
	assign w36085 = w36090 ^ w36050;
	assign w44881 = w36095 ^ w36098;
	assign w36048 = w36096 ^ w44881;
	assign w36004 = w36099 ^ w36048;
	assign w36086 = w47819 ^ w36004;
	assign w36084 = w36085 & w36086;
	assign w36082 = w36090 ^ w36084;
	assign w36003 = w36084 ^ w36048;
	assign w36002 = w36084 ^ w36101;
	assign w35997 = w36002 ^ w36098;
	assign w36008 = w36034 ^ w44881;
	assign w36092 = w36008 ^ w36033;
	assign w36083 = w36084 ^ w36092;
	assign w36089 = w36090 ^ w36092;
	assign w36088 = w36091 & w36089;
	assign w36087 = w36088 ^ w36050;
	assign w35999 = w36088 ^ w36100;
	assign w35995 = w35999 ^ w36035;
	assign w35998 = w47813 ^ w35995;
	assign w36075 = w35997 ^ w35998;
	assign w35996 = w36088 ^ w36044;
	assign w35994 = w47815 ^ w35995;
	assign w36081 = w36092 & w36082;
	assign w36079 = w36081 ^ w36089;
	assign w36078 = w36087 & w36079;
	assign w36043 = w36078 ^ w36053;
	assign w36077 = w36043 ^ w36045;
	assign w36001 = w36078 ^ w36102;
	assign w36074 = w36043 ^ w35996;
	assign w36069 = w36083 & w47820;
	assign w36068 = w36074 & w36104;
	assign w36067 = w36077 & w36116;
	assign w36066 = w36087 & w36106;
	assign w36010 = w36066 ^ w36067;
	assign w36065 = w36075 & w36107;
	assign w36060 = w36083 & w36115;
	assign w36059 = w36074 & w36119;
	assign w36026 = w36068 ^ w36059;
	assign w36058 = w36077 & w36112;
	assign w36028 = w36066 ^ w36058;
	assign w36057 = w36087 & w36113;
	assign w36056 = w36075 & w36118;
	assign w44882 = w36067 ^ w36068;
	assign w44884 = w36081 ^ w36099;
	assign w36040 = w47819 ^ w44884;
	assign w35993 = w36040 ^ w36001;
	assign w36000 = w36030 ^ w35993;
	assign w36076 = w35997 ^ w36000;
	assign w36072 = w35993 ^ w35994;
	assign w36064 = w36072 & w36105;
	assign w36025 = w36064 ^ w36067;
	assign w36022 = ~w36025;
	assign w36021 = w36064 ^ w36065;
	assign w36063 = w36076 & w36108;
	assign w36041 = w36059 ^ w36063;
	assign w36019 = ~w36041;
	assign w36018 = w36019 ^ w36057;
	assign w36055 = w36072 & w36120;
	assign w36054 = w36076 & w36117;
	assign w36020 = w36065 ^ w36054;
	assign w36016 = ~w36020;
	assign w43599 = w36055 ^ w36056;
	assign w36024 = w36028 ^ w43599;
	assign w36023 = w36019 ^ w36024;
	assign w36123 = w36022 ^ w36023;
	assign w36080 = w36040 ^ w36003;
	assign w36070 = w36080 & w36109;
	assign w36061 = w36080 & w36111;
	assign w36037 = w36061 ^ w43599;
	assign w36049 = w36064 ^ w44882;
	assign w36015 = w36060 ^ w36049;
	assign w36012 = ~w36015;
	assign w36009 = w36065 ^ w36049;
	assign w36073 = w44884 ^ w36051;
	assign w36071 = w36073 & w36110;
	assign w36062 = w36073 & w36114;
	assign w36038 = w36062 ^ w36037;
	assign w36042 = w36070 ^ w36038;
	assign w36047 = w36071 ^ w36042;
	assign w48443 = w44882 ^ w36047;
	assign w5972 = w48439 ^ w48443;
	assign w6098 = w48450 ^ w48443;
	assign w6108 = w5972 ^ w5973;
	assign w6110 = ~w6108;
	assign w6277 = w48453 ^ w48443;
	assign w5941 = w6278 ^ w6277;
	assign w48313 = w5941 ^ w5976;
	assign w47760 = w48313 ^ w4;
	assign w36122 = w36047 ^ w36021;
	assign w36011 = w36069 ^ w36042;
	assign w48442 = w36010 ^ w36011;
	assign w5963 = w48438 ^ w48442;
	assign w6081 = ~w5963;
	assign w6083 = w6081 ^ w5976;
	assign w6125 = w6124 ^ w48442;
	assign w48312 = w6126 ^ w6125;
	assign w47761 = w48312 ^ w3;
	assign w6240 = w48449 ^ w48442;
	assign w48446 = w36038 ^ w36009;
	assign w6027 = w48440 ^ w48446;
	assign w5938 = ~w6027;
	assign w6026 = w48446 ^ w48451;
	assign w6082 = w5938 ^ w48439;
	assign w48321 = w6083 ^ w6082;
	assign w47752 = w48321 ^ w12;
	assign w6092 = ~w6026;
	assign w6093 = w6092 ^ w48453;
	assign w6103 = w5938 ^ w48456;
	assign w6195 = w5533 ^ w48446;
	assign w6237 = w6027 ^ w48438;
	assign w6241 = w6026 ^ w48454;
	assign w5956 = w6241 ^ w6240;
	assign w48329 = w5956 ^ w5972;
	assign w48445 = ~w36122;
	assign w47744 = w48329 ^ w20;
	assign w44883 = w36069 ^ w36071;
	assign w36027 = w44883 ^ w36024;
	assign w36124 = w36026 ^ w36027;
	assign w36014 = w36018 ^ w44883;
	assign w36017 = w36056 ^ w36014;
	assign w36121 = w36016 ^ w36017;
	assign w6158 = w48454 ^ w36121;
	assign w36013 = w36037 ^ w36014;
	assign w48441 = w36012 ^ w36013;
	assign w5988 = w48441 ^ w48448;
	assign w6105 = ~w5988;
	assign w6094 = w5963 ^ w6105;
	assign w48328 = w6094 ^ w6093;
	assign w47745 = w48328 ^ w19;
	assign w6107 = w6105 ^ w48437;
	assign w6236 = w48437 ^ w48441;
	assign w5958 = w6237 ^ w6236;
	assign w48320 = w5958 ^ w5973;
	assign w47753 = w48320 ^ w11;
	assign w48444 = ~w36121;
	assign w44965 = w38105 ^ w38111;
	assign w38055 = w44965 ^ w38040;
	assign w38101 = w38063 ^ w38055;
	assign w38017 = w38049 ^ w44965;
	assign w38060 = w948 ^ w38017;
	assign w38095 = w38100 ^ w38060;
	assign w44966 = w38105 ^ w38108;
	assign w38058 = w38106 ^ w44966;
	assign w38014 = w38109 ^ w38058;
	assign w38096 = w944 ^ w38014;
	assign w38094 = w38095 & w38096;
	assign w38092 = w38100 ^ w38094;
	assign w38013 = w38094 ^ w38058;
	assign w38012 = w38094 ^ w38111;
	assign w38007 = w38012 ^ w38108;
	assign w38018 = w38044 ^ w44966;
	assign w38102 = w38018 ^ w38043;
	assign w38093 = w38094 ^ w38102;
	assign w38099 = w38100 ^ w38102;
	assign w38098 = w38101 & w38099;
	assign w38097 = w38098 ^ w38060;
	assign w38009 = w38098 ^ w38110;
	assign w38005 = w38009 ^ w38045;
	assign w38008 = w950 ^ w38005;
	assign w38085 = w38007 ^ w38008;
	assign w38006 = w38098 ^ w38054;
	assign w38004 = w948 ^ w38005;
	assign w38091 = w38102 & w38092;
	assign w38089 = w38091 ^ w38099;
	assign w38088 = w38097 & w38089;
	assign w38053 = w38088 ^ w38063;
	assign w38087 = w38053 ^ w38055;
	assign w38011 = w38088 ^ w38112;
	assign w38084 = w38053 ^ w38006;
	assign w38079 = w38093 & w943;
	assign w38078 = w38084 & w38114;
	assign w38077 = w38087 & w38126;
	assign w38076 = w38097 & w38116;
	assign w38020 = w38076 ^ w38077;
	assign w38075 = w38085 & w38117;
	assign w38070 = w38093 & w38125;
	assign w38069 = w38084 & w38129;
	assign w38036 = w38078 ^ w38069;
	assign w38068 = w38087 & w38122;
	assign w38038 = w38076 ^ w38068;
	assign w38067 = w38097 & w38123;
	assign w38066 = w38085 & w38128;
	assign w44967 = w38077 ^ w38078;
	assign w44969 = w38091 ^ w38109;
	assign w38050 = w944 ^ w44969;
	assign w38090 = w38050 ^ w38013;
	assign w38080 = w38090 & w38119;
	assign w38071 = w38090 & w38121;
	assign w38003 = w38050 ^ w38011;
	assign w38082 = w38003 ^ w38004;
	assign w38074 = w38082 & w38115;
	assign w38035 = w38074 ^ w38077;
	assign w38032 = ~w38035;
	assign w38031 = w38074 ^ w38075;
	assign w38065 = w38082 & w38130;
	assign w43604 = w38065 ^ w38066;
	assign w38034 = w38038 ^ w43604;
	assign w38047 = w38071 ^ w43604;
	assign w38059 = w38074 ^ w44967;
	assign w38025 = w38070 ^ w38059;
	assign w38022 = ~w38025;
	assign w38019 = w38075 ^ w38059;
	assign w38010 = w38040 ^ w38003;
	assign w38086 = w38007 ^ w38010;
	assign w38064 = w38086 & w38127;
	assign w38030 = w38075 ^ w38064;
	assign w38026 = ~w38030;
	assign w38073 = w38086 & w38118;
	assign w38051 = w38069 ^ w38073;
	assign w38029 = ~w38051;
	assign w38033 = w38029 ^ w38034;
	assign w38133 = w38032 ^ w38033;
	assign w48110 = ~w38133;
	assign w38028 = w38029 ^ w38067;
	assign w38083 = w44969 ^ w38061;
	assign w38081 = w38083 & w38120;
	assign w38072 = w38083 & w38124;
	assign w38048 = w38072 ^ w38047;
	assign w38052 = w38080 ^ w38048;
	assign w38057 = w38081 ^ w38052;
	assign w48113 = w44967 ^ w38057;
	assign w38132 = w38057 ^ w38031;
	assign w38021 = w38079 ^ w38052;
	assign w48112 = w38020 ^ w38021;
	assign w48116 = w38048 ^ w38019;
	assign w48115 = ~w38132;
	assign w44968 = w38079 ^ w38081;
	assign w38037 = w44968 ^ w38034;
	assign w38134 = w38036 ^ w38037;
	assign w48109 = ~w38134;
	assign w38024 = w38028 ^ w44968;
	assign w38027 = w38066 ^ w38024;
	assign w38131 = w38026 ^ w38027;
	assign w38023 = w38047 ^ w38024;
	assign w48111 = w38022 ^ w38023;
	assign w48114 = ~w38131;
	assign w44976 = w38373 ^ w38376;
	assign w38286 = w38312 ^ w44976;
	assign w38370 = w38286 ^ w38311;
	assign w38367 = w38368 ^ w38370;
	assign w38326 = w38374 ^ w44976;
	assign w38282 = w38377 ^ w38326;
	assign w38364 = w1709 ^ w38282;
	assign w44979 = w38373 ^ w38379;
	assign w38285 = w38317 ^ w44979;
	assign w38328 = w1713 ^ w38285;
	assign w38363 = w38368 ^ w38328;
	assign w38362 = w38363 & w38364;
	assign w38361 = w38362 ^ w38370;
	assign w38360 = w38368 ^ w38362;
	assign w38281 = w38362 ^ w38326;
	assign w38280 = w38362 ^ w38379;
	assign w38275 = w38280 ^ w38376;
	assign w38359 = w38370 & w38360;
	assign w38357 = w38359 ^ w38367;
	assign w38347 = w38361 & w1708;
	assign w38338 = w38361 & w38393;
	assign w44978 = w38359 ^ w38377;
	assign w38351 = w44978 ^ w38329;
	assign w38349 = w38351 & w38388;
	assign w38340 = w38351 & w38392;
	assign w38318 = w1709 ^ w44978;
	assign w38358 = w38318 ^ w38281;
	assign w38348 = w38358 & w38387;
	assign w38339 = w38358 & w38389;
	assign w38323 = w44979 ^ w38308;
	assign w38369 = w38331 ^ w38323;
	assign w38366 = w38369 & w38367;
	assign w38365 = w38366 ^ w38328;
	assign w38277 = w38366 ^ w38378;
	assign w38273 = w38277 ^ w38313;
	assign w38276 = w1715 ^ w38273;
	assign w38353 = w38275 ^ w38276;
	assign w38274 = w38366 ^ w38322;
	assign w38272 = w1713 ^ w38273;
	assign w38356 = w38365 & w38357;
	assign w38321 = w38356 ^ w38331;
	assign w38355 = w38321 ^ w38323;
	assign w38279 = w38356 ^ w38380;
	assign w38271 = w38318 ^ w38279;
	assign w38278 = w38308 ^ w38271;
	assign w38354 = w38275 ^ w38278;
	assign w38352 = w38321 ^ w38274;
	assign w38350 = w38271 ^ w38272;
	assign w38346 = w38352 & w38382;
	assign w38345 = w38355 & w38394;
	assign w38344 = w38365 & w38384;
	assign w38288 = w38344 ^ w38345;
	assign w38343 = w38353 & w38385;
	assign w38342 = w38350 & w38383;
	assign w38303 = w38342 ^ w38345;
	assign w38300 = ~w38303;
	assign w38299 = w38342 ^ w38343;
	assign w38341 = w38354 & w38386;
	assign w38337 = w38352 & w38397;
	assign w38319 = w38337 ^ w38341;
	assign w38304 = w38346 ^ w38337;
	assign w38297 = ~w38319;
	assign w38336 = w38355 & w38390;
	assign w38306 = w38344 ^ w38336;
	assign w38335 = w38365 & w38391;
	assign w38296 = w38297 ^ w38335;
	assign w38334 = w38353 & w38396;
	assign w38333 = w38350 & w38398;
	assign w38332 = w38354 & w38395;
	assign w38298 = w38343 ^ w38332;
	assign w38294 = ~w38298;
	assign w44977 = w38333 ^ w38334;
	assign w38315 = w38339 ^ w44977;
	assign w38316 = w38340 ^ w38315;
	assign w38320 = w38348 ^ w38316;
	assign w38325 = w38349 ^ w38320;
	assign w38400 = w38325 ^ w38299;
	assign w38289 = w38347 ^ w38320;
	assign w48048 = w38288 ^ w38289;
	assign w1750 = w1495 ^ w48048;
	assign w1782 = w1527 ^ w1750;
	assign w1814 = w1559 ^ w1782;
	assign w1846 = w1591 ^ w1814;
	assign w2045 = w1750 ^ w48112;
	assign w48051 = ~w38400;
	assign w1753 = w1498 ^ w48051;
	assign w1785 = w1530 ^ w1753;
	assign w1817 = w1562 ^ w1785;
	assign w1849 = w1594 ^ w1817;
	assign w988 = w1753 ^ w48115;
	assign w1020 = w1785 ^ w988;
	assign w1052 = w1817 ^ w1020;
	assign w1084 = w1849 ^ w1052;
	assign w38302 = w38306 ^ w44977;
	assign w38301 = w38297 ^ w38302;
	assign w38401 = w38300 ^ w38301;
	assign w48046 = ~w38401;
	assign w44980 = w38345 ^ w38346;
	assign w48049 = w44980 ^ w38325;
	assign w1751 = w1496 ^ w48049;
	assign w1783 = w1528 ^ w1751;
	assign w1815 = w1560 ^ w1783;
	assign w1847 = w1592 ^ w1815;
	assign w38176 = w1847 ^ w1849;
	assign w986 = w1751 ^ w48113;
	assign w1018 = w1783 ^ w986;
	assign w1050 = w1815 ^ w1018;
	assign w1082 = w1847 ^ w1050;
	assign w37908 = w1082 ^ w1084;
	assign w38327 = w38342 ^ w44980;
	assign w38293 = w38338 ^ w38327;
	assign w38290 = ~w38293;
	assign w38287 = w38343 ^ w38327;
	assign w48052 = w38316 ^ w38287;
	assign w1754 = w1499 ^ w48052;
	assign w1786 = w1531 ^ w1754;
	assign w1818 = w1563 ^ w1786;
	assign w1850 = w1595 ^ w1818;
	assign w989 = w1754 ^ w48116;
	assign w1021 = w1786 ^ w989;
	assign w1053 = w1818 ^ w1021;
	assign w1085 = w1850 ^ w1053;
	assign w37994 = w1082 ^ w1085;
	assign w38262 = w1847 ^ w1850;
	assign w44981 = w38347 ^ w38349;
	assign w38305 = w44981 ^ w38302;
	assign w38402 = w38304 ^ w38305;
	assign w48045 = ~w38402;
	assign w38292 = w38296 ^ w44981;
	assign w38295 = w38334 ^ w38292;
	assign w38399 = w38294 ^ w38295;
	assign w38291 = w38315 ^ w38292;
	assign w48047 = w38290 ^ w38291;
	assign w2044 = w1494 ^ w48047;
	assign w48050 = ~w38399;
	assign w1752 = w1497 ^ w48050;
	assign w1784 = w1529 ^ w1752;
	assign w1816 = w1561 ^ w1784;
	assign w1848 = w1593 ^ w1816;
	assign w987 = w1752 ^ w48114;
	assign w1019 = w1784 ^ w987;
	assign w1051 = w1816 ^ w1019;
	assign w1083 = w1848 ^ w1051;
	assign w37906 = w1083 ^ w1085;
	assign w37868 = w37908 ^ w37906;
	assign w37867 = w37908 ^ w1083;
	assign w38174 = w1848 ^ w1850;
	assign w38136 = w38176 ^ w38174;
	assign w38135 = w38176 ^ w1848;
	assign w44987 = w38641 ^ w38644;
	assign w38554 = w38580 ^ w44987;
	assign w38638 = w38554 ^ w38579;
	assign w38635 = w38636 ^ w38638;
	assign w38594 = w38642 ^ w44987;
	assign w38550 = w38645 ^ w38594;
	assign w38632 = w47891 ^ w38550;
	assign w44990 = w38641 ^ w38647;
	assign w38553 = w38585 ^ w44990;
	assign w38596 = w47887 ^ w38553;
	assign w38631 = w38636 ^ w38596;
	assign w38630 = w38631 & w38632;
	assign w38628 = w38636 ^ w38630;
	assign w38549 = w38630 ^ w38594;
	assign w38548 = w38630 ^ w38647;
	assign w38543 = w38548 ^ w38644;
	assign w38627 = w38638 & w38628;
	assign w38625 = w38627 ^ w38635;
	assign w44989 = w38627 ^ w38645;
	assign w38619 = w44989 ^ w38597;
	assign w38608 = w38619 & w38660;
	assign w38617 = w38619 & w38656;
	assign w38586 = w47891 ^ w44989;
	assign w38626 = w38586 ^ w38549;
	assign w38616 = w38626 & w38655;
	assign w38607 = w38626 & w38657;
	assign w38629 = w38630 ^ w38638;
	assign w38615 = w38629 & w47892;
	assign w38606 = w38629 & w38661;
	assign w38591 = w44990 ^ w38576;
	assign w38637 = w38599 ^ w38591;
	assign w38634 = w38637 & w38635;
	assign w38633 = w38634 ^ w38596;
	assign w38545 = w38634 ^ w38646;
	assign w38541 = w38545 ^ w38581;
	assign w38544 = w47885 ^ w38541;
	assign w38621 = w38543 ^ w38544;
	assign w38542 = w38634 ^ w38590;
	assign w38540 = w47887 ^ w38541;
	assign w38624 = w38633 & w38625;
	assign w38589 = w38624 ^ w38599;
	assign w38623 = w38589 ^ w38591;
	assign w38547 = w38624 ^ w38648;
	assign w38539 = w38586 ^ w38547;
	assign w38546 = w38576 ^ w38539;
	assign w38622 = w38543 ^ w38546;
	assign w38620 = w38589 ^ w38542;
	assign w38618 = w38539 ^ w38540;
	assign w38614 = w38620 & w38650;
	assign w38613 = w38623 & w38662;
	assign w38612 = w38633 & w38652;
	assign w38556 = w38612 ^ w38613;
	assign w38611 = w38621 & w38653;
	assign w38610 = w38618 & w38651;
	assign w38571 = w38610 ^ w38613;
	assign w38568 = ~w38571;
	assign w38567 = w38610 ^ w38611;
	assign w38609 = w38622 & w38654;
	assign w38605 = w38620 & w38665;
	assign w38587 = w38605 ^ w38609;
	assign w38572 = w38614 ^ w38605;
	assign w38565 = ~w38587;
	assign w38604 = w38623 & w38658;
	assign w38574 = w38612 ^ w38604;
	assign w38603 = w38633 & w38659;
	assign w38564 = w38565 ^ w38603;
	assign w38602 = w38621 & w38664;
	assign w38601 = w38618 & w38666;
	assign w38600 = w38622 & w38663;
	assign w38566 = w38611 ^ w38600;
	assign w38562 = ~w38566;
	assign w44988 = w38601 ^ w38602;
	assign w38583 = w38607 ^ w44988;
	assign w38584 = w38608 ^ w38583;
	assign w38588 = w38616 ^ w38584;
	assign w38557 = w38615 ^ w38588;
	assign w48494 = w38556 ^ w38557;
	assign w6008 = w48494 ^ w48507;
	assign w48424 = w5940 ^ w6008;
	assign w47649 = w48424 ^ w115;
	assign w6037 = w6008 ^ w6017;
	assign w38593 = w38617 ^ w38588;
	assign w38668 = w38593 ^ w38567;
	assign w6042 = w48501 ^ w38668;
	assign w48496 = ~w38668;
	assign w38570 = w38574 ^ w44988;
	assign w38569 = w38565 ^ w38570;
	assign w38669 = w38568 ^ w38569;
	assign w44991 = w38613 ^ w38614;
	assign w48495 = w44991 ^ w38593;
	assign w5968 = w48495 ^ w48500;
	assign w48433 = w5962 ^ w5968;
	assign w47640 = w48433 ^ w124;
	assign w6228 = ~w48495;
	assign w6229 = w48499 ^ w6228;
	assign w6039 = w48508 ^ w6228;
	assign w6063 = w5968 ^ w6014;
	assign w48425 = w6063 ^ w6062;
	assign w47648 = w48425 ^ w116;
	assign w38595 = w38610 ^ w44991;
	assign w38561 = w38606 ^ w38595;
	assign w38558 = ~w38561;
	assign w38555 = w38611 ^ w38595;
	assign w48497 = w38584 ^ w38555;
	assign w6033 = w48497 ^ w48501;
	assign w6022 = w48497 ^ w48509;
	assign w6036 = w6022 ^ w48500;
	assign w48409 = w6037 ^ w6036;
	assign w47664 = w48409 ^ w100;
	assign w6068 = w6033 ^ w48509;
	assign w44992 = w38615 ^ w38617;
	assign w38573 = w44992 ^ w38570;
	assign w38670 = w38572 ^ w38573;
	assign w38560 = w38564 ^ w44992;
	assign w38563 = w38602 ^ w38560;
	assign w38667 = w38562 ^ w38563;
	assign w38559 = w38583 ^ w38560;
	assign w48493 = w38558 ^ w38559;
	assign w5994 = w48493 ^ w48498;
	assign w6049 = w5994 ^ w6008;
	assign w6051 = ~w6049;
	assign w6061 = w5994 ^ w48506;
	assign w6266 = w6022 ^ w48493;
	assign w5946 = w6266 ^ w6265;
	assign w48408 = w5946 ^ w6014;
	assign w47665 = w48408 ^ w99;
	assign w45166 = ~w2043;
	assign w1525 = w1939 ^ w45166;
	assign w1557 = w1971 ^ w1525;
	assign w1589 = w2003 ^ w1557;
	assign w1749 = w45166 ^ w48046;
	assign w1780 = w1525 ^ w1749;
	assign w1812 = w1557 ^ w1780;
	assign w1844 = w1589 ^ w1812;
	assign w984 = w1749 ^ w48110;
	assign w1015 = w1780 ^ w984;
	assign w1047 = w1812 ^ w1015;
	assign w1079 = w1844 ^ w1047;
	assign w37995 = w1085 ^ w1079;
	assign w38173 = w1844 ^ w1846;
	assign w38254 = w38173 ^ w38262;
	assign w38252 = w38173 ^ w38136;
	assign w38263 = w1850 ^ w1844;
	assign w38441 = w1589 ^ w1591;
	assign w38443 = w1590 ^ w38441;
	assign w38519 = w1594 ^ w38443;
	assign w38516 = w1593 ^ w38443;
	assign w38522 = w38441 ^ w38530;
	assign w38458 = w1589 ^ w1590;
	assign w38526 = w38530 ^ w38458;
	assign w38520 = w38441 ^ w38404;
	assign w38531 = w1595 ^ w1589;
	assign w38515 = w38522 & w38526;
	assign w38447 = w38515 ^ w38444;
	assign w38512 = w38531 & w38516;
	assign w38446 = w38512 ^ w38442;
	assign w38509 = w38530 & w38519;
	assign w38445 = w38509 ^ w38443;
	assign w38451 = w38447 ^ w38445;
	assign w38456 = w1595 ^ w38451;
	assign w38417 = w38508 ^ w38509;
	assign w38464 = w38417 ^ w38418;
	assign w38463 = w38464 ^ w38446;
	assign w38507 = w38529 & w38520;
	assign w45167 = ~w2042;
	assign w1493 = w45167 ^ w47981;
	assign w1748 = w1493 ^ w48045;
	assign w983 = w1748 ^ w48109;
	assign w1938 = w216 ^ w45167;
	assign w1524 = w1938 ^ w1493;
	assign w1779 = w1524 ^ w1748;
	assign w1014 = w1779 ^ w983;
	assign w1970 = w184 ^ w1938;
	assign w2002 = w152 ^ w1970;
	assign w4178 = w2002 ^ w4179;
	assign w4104 = w2002 ^ w2008;
	assign w4175 = w4104 ^ w4099;
	assign w4182 = w4098 ^ w4104;
	assign w4180 = w4114 ^ w4182;
	assign w4185 = w2007 ^ w4104;
	assign w4181 = w2003 ^ w4185;
	assign w4184 = w2002 ^ w4059;
	assign w4171 = w4180 & w4178;
	assign w4121 = w4165 ^ w4171;
	assign w4163 = w4121 ^ w4112;
	assign w4170 = w4184 & w2002;
	assign w4168 = w4185 & w4181;
	assign w4162 = w4168 ^ w4119;
	assign w4167 = w4182 & w4175;
	assign w4159 = w4163 & w4162;
	assign w1556 = w1970 ^ w1524;
	assign w1588 = w2002 ^ w1556;
	assign w1811 = w1556 ^ w1779;
	assign w1843 = w1588 ^ w1811;
	assign w1046 = w1811 ^ w1014;
	assign w1078 = w1843 ^ w1046;
	assign w37912 = w1078 ^ w1084;
	assign w37989 = w37906 ^ w37912;
	assign w37992 = w1083 ^ w37912;
	assign w37988 = w1079 ^ w37992;
	assign w37991 = w1078 ^ w37867;
	assign w37977 = w37991 & w1078;
	assign w37975 = w37992 & w37988;
	assign w38253 = w1843 ^ w38254;
	assign w38180 = w1843 ^ w1849;
	assign w38257 = w38174 ^ w38180;
	assign w38260 = w1848 ^ w38180;
	assign w38256 = w1844 ^ w38260;
	assign w38259 = w1843 ^ w38135;
	assign w38245 = w38259 & w1843;
	assign w38243 = w38260 & w38256;
	assign w38521 = w1588 ^ w38522;
	assign w38448 = w1588 ^ w1594;
	assign w38518 = w38448 ^ w38443;
	assign w38525 = w38442 ^ w38448;
	assign w38523 = w38458 ^ w38525;
	assign w38528 = w1593 ^ w38448;
	assign w38524 = w1589 ^ w38528;
	assign w38527 = w1588 ^ w38403;
	assign w38514 = w38523 & w38521;
	assign w38465 = w38508 ^ w38514;
	assign w38506 = w38465 ^ w38456;
	assign w38513 = w38527 & w1588;
	assign w38511 = w38528 & w38524;
	assign w38505 = w38511 ^ w38463;
	assign w38510 = w38525 & w38518;
	assign w38502 = w38506 & w38505;
	assign w43704 = w4164 ^ w4170;
	assign w4075 = w4107 ^ w43704;
	assign w4118 = w2007 ^ w4075;
	assign w4154 = w4159 ^ w4118;
	assign w4113 = w43704 ^ w4098;
	assign w4160 = w4121 ^ w4113;
	assign w43705 = w4164 ^ w4167;
	assign w4116 = w4165 ^ w43705;
	assign w4072 = w4168 ^ w4116;
	assign w4155 = w2003 ^ w4072;
	assign w4153 = w4154 & w4155;
	assign w4071 = w4153 ^ w4116;
	assign w4070 = w4153 ^ w4170;
	assign w4065 = w4070 ^ w4167;
	assign w4151 = w4159 ^ w4153;
	assign w4076 = w4102 ^ w43705;
	assign w4161 = w4076 ^ w4101;
	assign w4152 = w4153 ^ w4161;
	assign w4150 = w4161 & w4151;
	assign w4138 = w4152 & w2002;
	assign w4129 = w4152 & w4184;
	assign w4158 = w4159 ^ w4161;
	assign w4148 = w4150 ^ w4158;
	assign w4157 = w4160 & w4158;
	assign w4067 = w4157 ^ w4169;
	assign w4063 = w4067 ^ w4103;
	assign w4066 = w2009 ^ w4063;
	assign w4144 = w4065 ^ w4066;
	assign w4064 = w4157 ^ w4112;
	assign w4062 = w2007 ^ w4063;
	assign w4134 = w4144 & w4176;
	assign w4125 = w4144 & w4187;
	assign w4156 = w4157 ^ w4118;
	assign w4147 = w4156 & w4148;
	assign w4069 = w4147 ^ w4171;
	assign w4135 = w4156 & w4175;
	assign w4126 = w4156 & w4182;
	assign w4111 = w4147 ^ w4121;
	assign w4146 = w4111 ^ w4113;
	assign w4143 = w4111 ^ w4064;
	assign w4137 = w4143 & w4173;
	assign w4136 = w4146 & w4185;
	assign w4078 = w4135 ^ w4136;
	assign w4128 = w4143 & w4188;
	assign w4127 = w4146 & w4181;
	assign w4094 = w4137 ^ w4128;
	assign w4096 = w4135 ^ w4127;
	assign w43706 = w4136 ^ w4137;
	assign w43708 = w4150 ^ w4168;
	assign w4142 = w43708 ^ w4119;
	assign w4140 = w4142 & w4179;
	assign w4131 = w4142 & w4183;
	assign w43707 = w4138 ^ w4140;
	assign w4108 = w2003 ^ w43708;
	assign w4061 = w4108 ^ w4069;
	assign w4068 = w4098 ^ w4061;
	assign w4149 = w4108 ^ w4071;
	assign w4139 = w4149 & w4178;
	assign w4130 = w4149 & w4180;
	assign w4141 = w4061 ^ w4062;
	assign w4133 = w4141 & w4174;
	assign w4145 = w4065 ^ w4068;
	assign w4132 = w4145 & w4177;
	assign w4124 = w4141 & w4189;
	assign w4123 = w4145 & w4186;
	assign w4122 = w4124 ^ w4125;
	assign w4105 = w4130 ^ w4122;
	assign w4106 = w4131 ^ w4105;
	assign w4109 = w4128 ^ w4132;
	assign w4110 = w4139 ^ w4106;
	assign w4079 = w4138 ^ w4110;
	assign w47952 = w4078 ^ w4079;
	assign w2037 = w123 ^ w47952;
	assign w1400 = w91 ^ w2037;
	assign w1432 = w59 ^ w1400;
	assign w1464 = w27 ^ w1432;
	assign w4117 = w4133 ^ w43706;
	assign w4077 = w4134 ^ w4117;
	assign w47956 = w4106 ^ w4077;
	assign w2041 = w127 ^ w47956;
	assign w1404 = w95 ^ w2041;
	assign w1436 = w63 ^ w1404;
	assign w1468 = w31 ^ w1436;
	assign w4083 = w4129 ^ w4117;
	assign w4080 = ~w4083;
	assign w4092 = w4096 ^ w4122;
	assign w4095 = w43707 ^ w4092;
	assign w4193 = w4094 ^ w4095;
	assign w47949 = ~w4193;
	assign w2034 = w120 ^ w47949;
	assign w1397 = w88 ^ w2034;
	assign w1429 = w56 ^ w1397;
	assign w1461 = w24 ^ w1429;
	assign w4115 = w4140 ^ w4110;
	assign w47953 = w43706 ^ w4115;
	assign w2038 = w124 ^ w47953;
	assign w1401 = w92 ^ w2038;
	assign w1433 = w60 ^ w1401;
	assign w1465 = w28 ^ w1433;
	assign w37458 = w1465 ^ w1468;
	assign w4089 = w4133 ^ w4134;
	assign w4191 = w4115 ^ w4089;
	assign w47955 = ~w4191;
	assign w2040 = w126 ^ w47955;
	assign w1403 = w94 ^ w2040;
	assign w1435 = w62 ^ w1403;
	assign w1467 = w30 ^ w1435;
	assign w37372 = w1465 ^ w1467;
	assign w37376 = w1461 ^ w1467;
	assign w4093 = w4133 ^ w4136;
	assign w4090 = ~w4093;
	assign w4087 = ~w4109;
	assign w4086 = w4087 ^ w4126;
	assign w4082 = w4086 ^ w43707;
	assign w4081 = w4105 ^ w4082;
	assign w47951 = w4080 ^ w4081;
	assign w2036 = w122 ^ w47951;
	assign w1399 = w90 ^ w2036;
	assign w1431 = w58 ^ w1399;
	assign w1463 = w26 ^ w1431;
	assign w37460 = w1463 ^ w1465;
	assign w37346 = w1464 ^ w1463;
	assign w37457 = w1468 ^ w1463;
	assign w4091 = w4087 ^ w4092;
	assign w4192 = w4090 ^ w4091;
	assign w47950 = ~w4192;
	assign w2035 = w121 ^ w47950;
	assign w1398 = w89 ^ w2035;
	assign w1430 = w57 ^ w1398;
	assign w1462 = w25 ^ w1430;
	assign w37369 = w1462 ^ w1464;
	assign w37371 = w1463 ^ w37369;
	assign w37447 = w1467 ^ w37371;
	assign w37446 = w37376 ^ w37371;
	assign w37450 = w37369 ^ w37458;
	assign w37449 = w1461 ^ w37450;
	assign w37386 = w1462 ^ w1463;
	assign w37454 = w37458 ^ w37386;
	assign w37459 = w1468 ^ w1462;
	assign w37443 = w37450 & w37454;
	assign w37375 = w37443 ^ w37372;
	assign w37437 = w37458 & w37447;
	assign w37373 = w37437 ^ w37371;
	assign w37379 = w37375 ^ w37373;
	assign w37384 = w1468 ^ w37379;
	assign w4088 = w4134 ^ w4123;
	assign w4084 = ~w4088;
	assign w4085 = w4125 ^ w4082;
	assign w4190 = w4084 ^ w4085;
	assign w47954 = ~w4190;
	assign w2039 = w125 ^ w47954;
	assign w1402 = w93 ^ w2039;
	assign w1434 = w61 ^ w1402;
	assign w1466 = w29 ^ w1434;
	assign w37444 = w1466 ^ w37371;
	assign w37370 = w1466 ^ w1468;
	assign w37445 = w37370 ^ w37460;
	assign w37453 = w37370 ^ w37376;
	assign w37451 = w37386 ^ w37453;
	assign w37456 = w1466 ^ w37376;
	assign w37452 = w1462 ^ w37456;
	assign w37332 = w37372 ^ w37370;
	assign w37448 = w37369 ^ w37332;
	assign w37331 = w37372 ^ w1466;
	assign w37455 = w1461 ^ w37331;
	assign w37442 = w37451 & w37449;
	assign w37441 = w37455 & w1461;
	assign w37440 = w37459 & w37444;
	assign w37374 = w37440 ^ w37370;
	assign w37439 = w37456 & w37452;
	assign w37438 = w37453 & w37446;
	assign w37436 = w37460 & w37445;
	assign w37393 = w37436 ^ w37442;
	assign w37434 = w37393 ^ w37384;
	assign w37345 = w37436 ^ w37437;
	assign w37392 = w37345 ^ w37346;
	assign w37391 = w37392 ^ w37374;
	assign w37433 = w37439 ^ w37391;
	assign w37435 = w37457 & w37448;
	assign w37430 = w37434 & w37433;
	assign w44936 = w37435 ^ w37441;
	assign w37347 = w37379 ^ w44936;
	assign w37390 = w1466 ^ w37347;
	assign w37425 = w37430 ^ w37390;
	assign w37385 = w44936 ^ w37370;
	assign w37431 = w37393 ^ w37385;
	assign w44937 = w37435 ^ w37438;
	assign w37388 = w37436 ^ w44937;
	assign w37344 = w37439 ^ w37388;
	assign w37426 = w1462 ^ w37344;
	assign w37424 = w37425 & w37426;
	assign w37422 = w37430 ^ w37424;
	assign w37343 = w37424 ^ w37388;
	assign w37342 = w37424 ^ w37441;
	assign w37337 = w37342 ^ w37438;
	assign w37348 = w37374 ^ w44937;
	assign w37432 = w37348 ^ w37373;
	assign w37423 = w37424 ^ w37432;
	assign w37429 = w37430 ^ w37432;
	assign w37428 = w37431 & w37429;
	assign w37427 = w37428 ^ w37390;
	assign w37339 = w37428 ^ w37440;
	assign w37335 = w37339 ^ w37375;
	assign w37338 = w1468 ^ w37335;
	assign w37415 = w37337 ^ w37338;
	assign w37336 = w37428 ^ w37384;
	assign w37334 = w1466 ^ w37335;
	assign w37421 = w37432 & w37422;
	assign w37419 = w37421 ^ w37429;
	assign w37418 = w37427 & w37419;
	assign w37383 = w37418 ^ w37393;
	assign w37417 = w37383 ^ w37385;
	assign w37341 = w37418 ^ w37442;
	assign w37414 = w37383 ^ w37336;
	assign w37409 = w37423 & w1461;
	assign w37408 = w37414 & w37444;
	assign w37407 = w37417 & w37456;
	assign w37406 = w37427 & w37446;
	assign w37350 = w37406 ^ w37407;
	assign w37405 = w37415 & w37447;
	assign w37400 = w37423 & w37455;
	assign w37399 = w37414 & w37459;
	assign w37366 = w37408 ^ w37399;
	assign w37398 = w37417 & w37452;
	assign w37368 = w37406 ^ w37398;
	assign w37397 = w37427 & w37453;
	assign w37396 = w37415 & w37458;
	assign w44939 = w37407 ^ w37408;
	assign w44941 = w37421 ^ w37439;
	assign w37413 = w44941 ^ w37391;
	assign w37402 = w37413 & w37454;
	assign w37411 = w37413 & w37450;
	assign w44940 = w37409 ^ w37411;
	assign w37380 = w1462 ^ w44941;
	assign w37420 = w37380 ^ w37343;
	assign w37333 = w37380 ^ w37341;
	assign w37340 = w37370 ^ w37333;
	assign w37416 = w37337 ^ w37340;
	assign w37412 = w37333 ^ w37334;
	assign w37410 = w37420 & w37449;
	assign w37404 = w37412 & w37445;
	assign w37389 = w37404 ^ w44939;
	assign w37365 = w37404 ^ w37407;
	assign w37362 = ~w37365;
	assign w37361 = w37404 ^ w37405;
	assign w37355 = w37400 ^ w37389;
	assign w37352 = ~w37355;
	assign w37349 = w37405 ^ w37389;
	assign w37403 = w37416 & w37448;
	assign w37381 = w37399 ^ w37403;
	assign w37359 = ~w37381;
	assign w37358 = w37359 ^ w37397;
	assign w37354 = w37358 ^ w44940;
	assign w37357 = w37396 ^ w37354;
	assign w37401 = w37420 & w37451;
	assign w37395 = w37412 & w37460;
	assign w37394 = w37416 & w37457;
	assign w37360 = w37405 ^ w37394;
	assign w37356 = ~w37360;
	assign w37461 = w37356 ^ w37357;
	assign w47962 = ~w37461;
	assign w1474 = w1888 ^ w47962;
	assign w1505 = w1919 ^ w1474;
	assign w1537 = w1951 ^ w1505;
	assign w1569 = w1983 ^ w1537;
	assign w44938 = w37395 ^ w37396;
	assign w37364 = w37368 ^ w44938;
	assign w37367 = w44940 ^ w37364;
	assign w37464 = w37366 ^ w37367;
	assign w47957 = ~w37464;
	assign w1469 = w1883 ^ w47957;
	assign w1500 = w1914 ^ w1469;
	assign w1532 = w1946 ^ w1500;
	assign w1564 = w1978 ^ w1532;
	assign w37363 = w37359 ^ w37364;
	assign w37463 = w37362 ^ w37363;
	assign w47958 = ~w37463;
	assign w1470 = w1884 ^ w47958;
	assign w1501 = w1915 ^ w1470;
	assign w1533 = w1947 ^ w1501;
	assign w1565 = w1979 ^ w1533;
	assign w37377 = w37401 ^ w44938;
	assign w37378 = w37402 ^ w37377;
	assign w37382 = w37410 ^ w37378;
	assign w37387 = w37411 ^ w37382;
	assign w47961 = w44939 ^ w37387;
	assign w1473 = w1887 ^ w47961;
	assign w1504 = w1918 ^ w1473;
	assign w1536 = w1950 ^ w1504;
	assign w1568 = w1982 ^ w1536;
	assign w37462 = w37387 ^ w37361;
	assign w37353 = w37377 ^ w37354;
	assign w47959 = w37352 ^ w37353;
	assign w1471 = w1885 ^ w47959;
	assign w1502 = w1916 ^ w1471;
	assign w1534 = w1948 ^ w1502;
	assign w1566 = w1980 ^ w1534;
	assign w37252 = w1565 ^ w1566;
	assign w37326 = w1566 ^ w1568;
	assign w37351 = w37409 ^ w37382;
	assign w47960 = w37350 ^ w37351;
	assign w1472 = w1886 ^ w47960;
	assign w1503 = w1917 ^ w1472;
	assign w1535 = w1949 ^ w1503;
	assign w1567 = w1981 ^ w1535;
	assign w37235 = w1565 ^ w1567;
	assign w37237 = w1566 ^ w37235;
	assign w37310 = w1569 ^ w37237;
	assign w37212 = w1567 ^ w1566;
	assign w47964 = w37378 ^ w37349;
	assign w1476 = w1890 ^ w47964;
	assign w1507 = w1921 ^ w1476;
	assign w1539 = w1953 ^ w1507;
	assign w1571 = w1985 ^ w1539;
	assign w37236 = w1569 ^ w1571;
	assign w37311 = w37236 ^ w37326;
	assign w37324 = w1568 ^ w1571;
	assign w37320 = w37324 ^ w37252;
	assign w37316 = w37235 ^ w37324;
	assign w37315 = w1564 ^ w37316;
	assign w37325 = w1571 ^ w1565;
	assign w37323 = w1571 ^ w1566;
	assign w37309 = w37316 & w37320;
	assign w37306 = w37325 & w37310;
	assign w37240 = w37306 ^ w37236;
	assign w37302 = w37326 & w37311;
	assign w47963 = ~w37462;
	assign w1475 = w1889 ^ w47963;
	assign w1506 = w1920 ^ w1475;
	assign w1538 = w1952 ^ w1506;
	assign w1570 = w1984 ^ w1538;
	assign w37313 = w1570 ^ w37237;
	assign w37238 = w1568 ^ w1570;
	assign w37241 = w37309 ^ w37238;
	assign w37242 = w1564 ^ w1570;
	assign w37312 = w37242 ^ w37237;
	assign w37319 = w37236 ^ w37242;
	assign w37317 = w37252 ^ w37319;
	assign w37322 = w1569 ^ w37242;
	assign w37318 = w1565 ^ w37322;
	assign w37198 = w37238 ^ w37236;
	assign w37314 = w37235 ^ w37198;
	assign w37197 = w37238 ^ w1569;
	assign w37321 = w1564 ^ w37197;
	assign w37308 = w37317 & w37315;
	assign w37259 = w37302 ^ w37308;
	assign w37307 = w37321 & w1564;
	assign w37305 = w37322 & w37318;
	assign w37304 = w37319 & w37312;
	assign w37303 = w37324 & w37313;
	assign w37239 = w37303 ^ w37237;
	assign w37245 = w37241 ^ w37239;
	assign w37250 = w1571 ^ w37245;
	assign w37300 = w37259 ^ w37250;
	assign w37211 = w37302 ^ w37303;
	assign w37258 = w37211 ^ w37212;
	assign w37257 = w37258 ^ w37240;
	assign w37299 = w37305 ^ w37257;
	assign w37301 = w37323 & w37314;
	assign w37296 = w37300 & w37299;
	assign w44931 = w37301 ^ w37307;
	assign w37251 = w44931 ^ w37236;
	assign w37297 = w37259 ^ w37251;
	assign w37213 = w37245 ^ w44931;
	assign w37256 = w1569 ^ w37213;
	assign w37291 = w37296 ^ w37256;
	assign w44932 = w37301 ^ w37304;
	assign w37254 = w37302 ^ w44932;
	assign w37210 = w37305 ^ w37254;
	assign w37292 = w1565 ^ w37210;
	assign w37290 = w37291 & w37292;
	assign w37288 = w37296 ^ w37290;
	assign w37209 = w37290 ^ w37254;
	assign w37208 = w37290 ^ w37307;
	assign w37203 = w37208 ^ w37304;
	assign w37214 = w37240 ^ w44932;
	assign w37298 = w37214 ^ w37239;
	assign w37289 = w37290 ^ w37298;
	assign w37295 = w37296 ^ w37298;
	assign w37294 = w37297 & w37295;
	assign w37293 = w37294 ^ w37256;
	assign w37205 = w37294 ^ w37306;
	assign w37201 = w37205 ^ w37241;
	assign w37204 = w1571 ^ w37201;
	assign w37281 = w37203 ^ w37204;
	assign w37202 = w37294 ^ w37250;
	assign w37200 = w1569 ^ w37201;
	assign w37287 = w37298 & w37288;
	assign w37285 = w37287 ^ w37295;
	assign w37284 = w37293 & w37285;
	assign w37249 = w37284 ^ w37259;
	assign w37283 = w37249 ^ w37251;
	assign w37207 = w37284 ^ w37308;
	assign w37280 = w37249 ^ w37202;
	assign w37275 = w37289 & w1564;
	assign w37274 = w37280 & w37310;
	assign w37273 = w37283 & w37322;
	assign w37272 = w37293 & w37312;
	assign w37216 = w37272 ^ w37273;
	assign w37271 = w37281 & w37313;
	assign w37266 = w37289 & w37321;
	assign w37265 = w37280 & w37325;
	assign w37232 = w37274 ^ w37265;
	assign w37264 = w37283 & w37318;
	assign w37234 = w37272 ^ w37264;
	assign w37263 = w37293 & w37319;
	assign w37262 = w37281 & w37324;
	assign w44933 = w37273 ^ w37274;
	assign w44935 = w37287 ^ w37305;
	assign w37246 = w1565 ^ w44935;
	assign w37199 = w37246 ^ w37207;
	assign w37206 = w37236 ^ w37199;
	assign w37282 = w37203 ^ w37206;
	assign w37269 = w37282 & w37314;
	assign w37247 = w37265 ^ w37269;
	assign w37225 = ~w37247;
	assign w37278 = w37199 ^ w37200;
	assign w37270 = w37278 & w37311;
	assign w37227 = w37270 ^ w37271;
	assign w37231 = w37270 ^ w37273;
	assign w37228 = ~w37231;
	assign w37224 = w37225 ^ w37263;
	assign w37261 = w37278 & w37326;
	assign w37260 = w37282 & w37323;
	assign w37226 = w37271 ^ w37260;
	assign w37222 = ~w37226;
	assign w43602 = w37261 ^ w37262;
	assign w37230 = w37234 ^ w43602;
	assign w37229 = w37225 ^ w37230;
	assign w37329 = w37228 ^ w37229;
	assign w47990 = ~w37329;
	assign w1597 = w2011 ^ w47990;
	assign w1629 = w1374 ^ w1597;
	assign w1661 = w1406 ^ w1629;
	assign w1693 = w1438 ^ w1661;
	assign w37286 = w37246 ^ w37209;
	assign w37276 = w37286 & w37315;
	assign w37267 = w37286 & w37317;
	assign w37243 = w37267 ^ w43602;
	assign w37255 = w37270 ^ w44933;
	assign w37221 = w37266 ^ w37255;
	assign w37218 = ~w37221;
	assign w37215 = w37271 ^ w37255;
	assign w37279 = w44935 ^ w37257;
	assign w37277 = w37279 & w37316;
	assign w37268 = w37279 & w37320;
	assign w37244 = w37268 ^ w37243;
	assign w37248 = w37276 ^ w37244;
	assign w37253 = w37277 ^ w37248;
	assign w47993 = w44933 ^ w37253;
	assign w1600 = w2014 ^ w47993;
	assign w1632 = w1377 ^ w1600;
	assign w1664 = w1409 ^ w1632;
	assign w1696 = w1441 ^ w1664;
	assign w37328 = w37253 ^ w37227;
	assign w37217 = w37275 ^ w37248;
	assign w47992 = w37216 ^ w37217;
	assign w1599 = w2013 ^ w47992;
	assign w1631 = w1376 ^ w1599;
	assign w1663 = w1408 ^ w1631;
	assign w1695 = w1440 ^ w1663;
	assign w23165 = w1693 ^ w1695;
	assign w47996 = w37244 ^ w37215;
	assign w1603 = w2017 ^ w47996;
	assign w1635 = w1380 ^ w1603;
	assign w1667 = w1412 ^ w1635;
	assign w1699 = w1444 ^ w1667;
	assign w23254 = w1696 ^ w1699;
	assign w23246 = w23165 ^ w23254;
	assign w23255 = w1699 ^ w1693;
	assign w47995 = ~w37328;
	assign w1602 = w2016 ^ w47995;
	assign w1634 = w1379 ^ w1602;
	assign w1666 = w1411 ^ w1634;
	assign w1698 = w1443 ^ w1666;
	assign w23168 = w1696 ^ w1698;
	assign w44934 = w37275 ^ w37277;
	assign w37233 = w44934 ^ w37230;
	assign w37330 = w37232 ^ w37233;
	assign w47989 = ~w37330;
	assign w1596 = w2010 ^ w47989;
	assign w1628 = w1373 ^ w1596;
	assign w1660 = w1405 ^ w1628;
	assign w1692 = w1437 ^ w1660;
	assign w23245 = w1692 ^ w23246;
	assign w23172 = w1692 ^ w1698;
	assign w37220 = w37224 ^ w44934;
	assign w37223 = w37262 ^ w37220;
	assign w37327 = w37222 ^ w37223;
	assign w37219 = w37243 ^ w37220;
	assign w47991 = w37218 ^ w37219;
	assign w1598 = w2012 ^ w47991;
	assign w1630 = w1375 ^ w1598;
	assign w1662 = w1407 ^ w1630;
	assign w1694 = w1439 ^ w1662;
	assign w23167 = w1694 ^ w23165;
	assign w23243 = w1698 ^ w23167;
	assign w23242 = w23172 ^ w23167;
	assign w23182 = w1693 ^ w1694;
	assign w23250 = w23254 ^ w23182;
	assign w23256 = w1694 ^ w1696;
	assign w23142 = w1695 ^ w1694;
	assign w23253 = w1699 ^ w1694;
	assign w23239 = w23246 & w23250;
	assign w23171 = w23239 ^ w23168;
	assign w23233 = w23254 & w23243;
	assign w23169 = w23233 ^ w23167;
	assign w23175 = w23171 ^ w23169;
	assign w23180 = w1699 ^ w23175;
	assign w47994 = ~w37327;
	assign w1601 = w2015 ^ w47994;
	assign w1633 = w1378 ^ w1601;
	assign w1665 = w1410 ^ w1633;
	assign w1697 = w1442 ^ w1665;
	assign w23240 = w1697 ^ w23167;
	assign w23166 = w1697 ^ w1699;
	assign w23241 = w23166 ^ w23256;
	assign w23249 = w23166 ^ w23172;
	assign w23247 = w23182 ^ w23249;
	assign w23252 = w1697 ^ w23172;
	assign w23248 = w1693 ^ w23252;
	assign w23128 = w23168 ^ w23166;
	assign w23244 = w23165 ^ w23128;
	assign w23127 = w23168 ^ w1697;
	assign w23251 = w1692 ^ w23127;
	assign w23238 = w23247 & w23245;
	assign w23237 = w23251 & w1692;
	assign w23236 = w23255 & w23240;
	assign w23170 = w23236 ^ w23166;
	assign w23235 = w23252 & w23248;
	assign w23234 = w23249 & w23242;
	assign w23232 = w23256 & w23241;
	assign w23189 = w23232 ^ w23238;
	assign w23230 = w23189 ^ w23180;
	assign w23141 = w23232 ^ w23233;
	assign w23188 = w23141 ^ w23142;
	assign w23187 = w23188 ^ w23170;
	assign w23229 = w23235 ^ w23187;
	assign w23231 = w23253 & w23244;
	assign w23226 = w23230 & w23229;
	assign w44340 = w23231 ^ w23234;
	assign w23144 = w23170 ^ w44340;
	assign w23228 = w23144 ^ w23169;
	assign w23225 = w23226 ^ w23228;
	assign w23184 = w23232 ^ w44340;
	assign w23140 = w23235 ^ w23184;
	assign w23222 = w1693 ^ w23140;
	assign w44343 = w23231 ^ w23237;
	assign w23143 = w23175 ^ w44343;
	assign w23186 = w1697 ^ w23143;
	assign w23221 = w23226 ^ w23186;
	assign w23220 = w23221 & w23222;
	assign w23219 = w23220 ^ w23228;
	assign w23218 = w23226 ^ w23220;
	assign w23139 = w23220 ^ w23184;
	assign w23138 = w23220 ^ w23237;
	assign w23133 = w23138 ^ w23234;
	assign w23217 = w23228 & w23218;
	assign w23215 = w23217 ^ w23225;
	assign w23205 = w23219 & w1692;
	assign w23196 = w23219 & w23251;
	assign w44342 = w23217 ^ w23235;
	assign w23209 = w44342 ^ w23187;
	assign w23207 = w23209 & w23246;
	assign w23198 = w23209 & w23250;
	assign w23176 = w1693 ^ w44342;
	assign w23216 = w23176 ^ w23139;
	assign w23206 = w23216 & w23245;
	assign w23197 = w23216 & w23247;
	assign w23181 = w44343 ^ w23166;
	assign w23227 = w23189 ^ w23181;
	assign w23224 = w23227 & w23225;
	assign w23223 = w23224 ^ w23186;
	assign w23135 = w23224 ^ w23236;
	assign w23131 = w23135 ^ w23171;
	assign w23134 = w1699 ^ w23131;
	assign w23211 = w23133 ^ w23134;
	assign w23132 = w23224 ^ w23180;
	assign w23130 = w1697 ^ w23131;
	assign w23214 = w23223 & w23215;
	assign w23179 = w23214 ^ w23189;
	assign w23213 = w23179 ^ w23181;
	assign w23137 = w23214 ^ w23238;
	assign w23129 = w23176 ^ w23137;
	assign w23136 = w23166 ^ w23129;
	assign w23212 = w23133 ^ w23136;
	assign w23210 = w23179 ^ w23132;
	assign w23208 = w23129 ^ w23130;
	assign w23204 = w23210 & w23240;
	assign w23203 = w23213 & w23252;
	assign w23202 = w23223 & w23242;
	assign w23146 = w23202 ^ w23203;
	assign w23201 = w23211 & w23243;
	assign w23200 = w23208 & w23241;
	assign w23161 = w23200 ^ w23203;
	assign w23158 = ~w23161;
	assign w23157 = w23200 ^ w23201;
	assign w23199 = w23212 & w23244;
	assign w23195 = w23210 & w23255;
	assign w23177 = w23195 ^ w23199;
	assign w23162 = w23204 ^ w23195;
	assign w23155 = ~w23177;
	assign w23194 = w23213 & w23248;
	assign w23164 = w23202 ^ w23194;
	assign w23193 = w23223 & w23249;
	assign w23154 = w23155 ^ w23193;
	assign w23192 = w23211 & w23254;
	assign w23191 = w23208 & w23256;
	assign w23190 = w23212 & w23253;
	assign w23156 = w23201 ^ w23190;
	assign w23152 = ~w23156;
	assign w44341 = w23191 ^ w23192;
	assign w23173 = w23197 ^ w44341;
	assign w23174 = w23198 ^ w23173;
	assign w23178 = w23206 ^ w23174;
	assign w23183 = w23207 ^ w23178;
	assign w23258 = w23183 ^ w23157;
	assign w23147 = w23205 ^ w23178;
	assign w48032 = w23146 ^ w23147;
	assign w1735 = w1480 ^ w48032;
	assign w1766 = w1511 ^ w1735;
	assign w1798 = w1543 ^ w1766;
	assign w1830 = w1575 ^ w1798;
	assign w48035 = ~w23258;
	assign w1738 = w1483 ^ w48035;
	assign w1769 = w1514 ^ w1738;
	assign w1801 = w1546 ^ w1769;
	assign w1833 = w1578 ^ w1801;
	assign w23160 = w23164 ^ w44341;
	assign w23159 = w23155 ^ w23160;
	assign w23259 = w23158 ^ w23159;
	assign w48030 = ~w23259;
	assign w1733 = w1478 ^ w48030;
	assign w1764 = w1509 ^ w1733;
	assign w1796 = w1541 ^ w1764;
	assign w1828 = w1573 ^ w1796;
	assign w23031 = w1828 ^ w1830;
	assign w44344 = w23203 ^ w23204;
	assign w48033 = w44344 ^ w23183;
	assign w1736 = w1481 ^ w48033;
	assign w1767 = w1512 ^ w1736;
	assign w1799 = w1544 ^ w1767;
	assign w1831 = w1576 ^ w1799;
	assign w23034 = w1831 ^ w1833;
	assign w23185 = w23200 ^ w44344;
	assign w23151 = w23196 ^ w23185;
	assign w23148 = ~w23151;
	assign w23145 = w23201 ^ w23185;
	assign w48036 = w23174 ^ w23145;
	assign w1739 = w1484 ^ w48036;
	assign w1770 = w1515 ^ w1739;
	assign w1802 = w1547 ^ w1770;
	assign w1834 = w1579 ^ w1802;
	assign w23120 = w1831 ^ w1834;
	assign w23112 = w23031 ^ w23120;
	assign w23121 = w1834 ^ w1828;
	assign w44345 = w23205 ^ w23207;
	assign w23163 = w44345 ^ w23160;
	assign w23260 = w23162 ^ w23163;
	assign w48029 = ~w23260;
	assign w1732 = w1477 ^ w48029;
	assign w1763 = w1508 ^ w1732;
	assign w1795 = w1540 ^ w1763;
	assign w1827 = w1572 ^ w1795;
	assign w23038 = w1827 ^ w1833;
	assign w23111 = w1827 ^ w23112;
	assign w23150 = w23154 ^ w44345;
	assign w23153 = w23192 ^ w23150;
	assign w23257 = w23152 ^ w23153;
	assign w23149 = w23173 ^ w23150;
	assign w48031 = w23148 ^ w23149;
	assign w1734 = w1479 ^ w48031;
	assign w1765 = w1510 ^ w1734;
	assign w1797 = w1542 ^ w1765;
	assign w1829 = w1574 ^ w1797;
	assign w23033 = w1829 ^ w23031;
	assign w23109 = w1833 ^ w23033;
	assign w23108 = w23038 ^ w23033;
	assign w23048 = w1828 ^ w1829;
	assign w23116 = w23120 ^ w23048;
	assign w23122 = w1829 ^ w1831;
	assign w23008 = w1830 ^ w1829;
	assign w23119 = w1834 ^ w1829;
	assign w23105 = w23112 & w23116;
	assign w23037 = w23105 ^ w23034;
	assign w23099 = w23120 & w23109;
	assign w23035 = w23099 ^ w23033;
	assign w23041 = w23037 ^ w23035;
	assign w23046 = w1834 ^ w23041;
	assign w48034 = ~w23257;
	assign w1737 = w1482 ^ w48034;
	assign w1768 = w1513 ^ w1737;
	assign w1800 = w1545 ^ w1768;
	assign w1832 = w1577 ^ w1800;
	assign w23106 = w1832 ^ w23033;
	assign w23032 = w1832 ^ w1834;
	assign w23107 = w23032 ^ w23122;
	assign w23115 = w23032 ^ w23038;
	assign w23113 = w23048 ^ w23115;
	assign w23118 = w1832 ^ w23038;
	assign w23114 = w1828 ^ w23118;
	assign w22994 = w23034 ^ w23032;
	assign w23110 = w23031 ^ w22994;
	assign w22993 = w23034 ^ w1832;
	assign w23117 = w1827 ^ w22993;
	assign w23104 = w23113 & w23111;
	assign w23103 = w23117 & w1827;
	assign w23102 = w23121 & w23106;
	assign w23036 = w23102 ^ w23032;
	assign w23101 = w23118 & w23114;
	assign w23100 = w23115 & w23108;
	assign w23098 = w23122 & w23107;
	assign w23055 = w23098 ^ w23104;
	assign w23096 = w23055 ^ w23046;
	assign w23007 = w23098 ^ w23099;
	assign w23054 = w23007 ^ w23008;
	assign w23053 = w23054 ^ w23036;
	assign w23095 = w23101 ^ w23053;
	assign w23097 = w23119 & w23110;
	assign w23092 = w23096 & w23095;
	assign w44334 = w23097 ^ w23103;
	assign w23009 = w23041 ^ w44334;
	assign w23052 = w1832 ^ w23009;
	assign w23087 = w23092 ^ w23052;
	assign w23047 = w44334 ^ w23032;
	assign w23093 = w23055 ^ w23047;
	assign w44335 = w23097 ^ w23100;
	assign w23050 = w23098 ^ w44335;
	assign w23006 = w23101 ^ w23050;
	assign w23088 = w1828 ^ w23006;
	assign w23086 = w23087 & w23088;
	assign w23084 = w23092 ^ w23086;
	assign w23005 = w23086 ^ w23050;
	assign w23004 = w23086 ^ w23103;
	assign w22999 = w23004 ^ w23100;
	assign w23010 = w23036 ^ w44335;
	assign w23094 = w23010 ^ w23035;
	assign w23085 = w23086 ^ w23094;
	assign w23091 = w23092 ^ w23094;
	assign w23090 = w23093 & w23091;
	assign w23089 = w23090 ^ w23052;
	assign w23001 = w23090 ^ w23102;
	assign w22997 = w23001 ^ w23037;
	assign w23000 = w1834 ^ w22997;
	assign w23077 = w22999 ^ w23000;
	assign w22998 = w23090 ^ w23046;
	assign w22996 = w1832 ^ w22997;
	assign w23083 = w23094 & w23084;
	assign w23081 = w23083 ^ w23091;
	assign w23080 = w23089 & w23081;
	assign w23045 = w23080 ^ w23055;
	assign w23079 = w23045 ^ w23047;
	assign w23003 = w23080 ^ w23104;
	assign w23076 = w23045 ^ w22998;
	assign w23071 = w23085 & w1827;
	assign w23070 = w23076 & w23106;
	assign w23069 = w23079 & w23118;
	assign w23068 = w23089 & w23108;
	assign w23012 = w23068 ^ w23069;
	assign w23067 = w23077 & w23109;
	assign w23062 = w23085 & w23117;
	assign w23061 = w23076 & w23121;
	assign w23028 = w23070 ^ w23061;
	assign w23060 = w23079 & w23114;
	assign w23030 = w23068 ^ w23060;
	assign w23059 = w23089 & w23115;
	assign w23058 = w23077 & w23120;
	assign w44337 = w23069 ^ w23070;
	assign w44339 = w23083 ^ w23101;
	assign w23075 = w44339 ^ w23053;
	assign w23064 = w23075 & w23116;
	assign w23073 = w23075 & w23112;
	assign w44338 = w23071 ^ w23073;
	assign w23042 = w1828 ^ w44339;
	assign w23082 = w23042 ^ w23005;
	assign w22995 = w23042 ^ w23003;
	assign w23002 = w23032 ^ w22995;
	assign w23078 = w22999 ^ w23002;
	assign w23074 = w22995 ^ w22996;
	assign w23072 = w23082 & w23111;
	assign w23066 = w23074 & w23107;
	assign w23051 = w23066 ^ w44337;
	assign w23027 = w23066 ^ w23069;
	assign w23024 = ~w23027;
	assign w23023 = w23066 ^ w23067;
	assign w23017 = w23062 ^ w23051;
	assign w23014 = ~w23017;
	assign w23011 = w23067 ^ w23051;
	assign w23065 = w23078 & w23110;
	assign w23043 = w23061 ^ w23065;
	assign w23021 = ~w23043;
	assign w23020 = w23021 ^ w23059;
	assign w23016 = w23020 ^ w44338;
	assign w23019 = w23058 ^ w23016;
	assign w23063 = w23082 & w23113;
	assign w23057 = w23074 & w23122;
	assign w23056 = w23078 & w23119;
	assign w23022 = w23067 ^ w23056;
	assign w23018 = ~w23022;
	assign w23123 = w23018 ^ w23019;
	assign w48066 = ~w23123;
	assign w1864 = w1609 ^ w48066;
	assign w876 = w1641 ^ w1864;
	assign w908 = w1673 ^ w876;
	assign w940 = w1705 ^ w908;
	assign w44336 = w23057 ^ w23058;
	assign w23039 = w23063 ^ w44336;
	assign w23015 = w23039 ^ w23016;
	assign w48063 = w23014 ^ w23015;
	assign w1861 = w1606 ^ w48063;
	assign w873 = w1638 ^ w1861;
	assign w905 = w1670 ^ w873;
	assign w23040 = w23064 ^ w23039;
	assign w48068 = w23040 ^ w23011;
	assign w1866 = w1611 ^ w48068;
	assign w878 = w1643 ^ w1866;
	assign w910 = w1675 ^ w878;
	assign w23044 = w23072 ^ w23040;
	assign w23013 = w23071 ^ w23044;
	assign w48064 = w23012 ^ w23013;
	assign w1862 = w1607 ^ w48064;
	assign w874 = w1639 ^ w1862;
	assign w906 = w1671 ^ w874;
	assign w938 = w1703 ^ w906;
	assign w942 = w1707 ^ w910;
	assign w23049 = w23073 ^ w23044;
	assign w23124 = w23049 ^ w23023;
	assign w48067 = ~w23124;
	assign w1865 = w1610 ^ w48067;
	assign w877 = w1642 ^ w1865;
	assign w909 = w1674 ^ w877;
	assign w941 = w1706 ^ w909;
	assign w937 = w1702 ^ w905;
	assign w35226 = w940 ^ w942;
	assign w35202 = w938 ^ w937;
	assign w35313 = w942 ^ w937;
	assign w48065 = w44337 ^ w23049;
	assign w1863 = w1608 ^ w48065;
	assign w875 = w1640 ^ w1863;
	assign w907 = w1672 ^ w875;
	assign w939 = w1704 ^ w907;
	assign w35228 = w939 ^ w941;
	assign w35314 = w939 ^ w942;
	assign w35316 = w937 ^ w939;
	assign w35301 = w35226 ^ w35316;
	assign w35188 = w35228 ^ w35226;
	assign w35187 = w35228 ^ w940;
	assign w35292 = w35316 & w35301;
	assign w23026 = w23030 ^ w44336;
	assign w23029 = w44338 ^ w23026;
	assign w23126 = w23028 ^ w23029;
	assign w23025 = w23021 ^ w23026;
	assign w23125 = w23024 ^ w23025;
	assign w48061 = ~w23126;
	assign w1859 = w1604 ^ w48061;
	assign w871 = w1636 ^ w1859;
	assign w903 = w1668 ^ w871;
	assign w48062 = ~w23125;
	assign w1860 = w1605 ^ w48062;
	assign w872 = w1637 ^ w1860;
	assign w904 = w1669 ^ w872;
	assign w936 = w1701 ^ w904;
	assign w935 = w1700 ^ w903;
	assign w35225 = w936 ^ w938;
	assign w35227 = w937 ^ w35225;
	assign w35303 = w941 ^ w35227;
	assign w35300 = w940 ^ w35227;
	assign w35232 = w935 ^ w941;
	assign w35302 = w35232 ^ w35227;
	assign w35309 = w35226 ^ w35232;
	assign w35306 = w35225 ^ w35314;
	assign w35305 = w935 ^ w35306;
	assign w35242 = w936 ^ w937;
	assign w35307 = w35242 ^ w35309;
	assign w35310 = w35314 ^ w35242;
	assign w35312 = w940 ^ w35232;
	assign w35308 = w936 ^ w35312;
	assign w35304 = w35225 ^ w35188;
	assign w35311 = w935 ^ w35187;
	assign w35315 = w942 ^ w936;
	assign w35299 = w35306 & w35310;
	assign w35231 = w35299 ^ w35228;
	assign w35298 = w35307 & w35305;
	assign w35249 = w35292 ^ w35298;
	assign w35297 = w35311 & w935;
	assign w35296 = w35315 & w35300;
	assign w35230 = w35296 ^ w35226;
	assign w35295 = w35312 & w35308;
	assign w35294 = w35309 & w35302;
	assign w35293 = w35314 & w35303;
	assign w35229 = w35293 ^ w35227;
	assign w35235 = w35231 ^ w35229;
	assign w35240 = w942 ^ w35235;
	assign w35290 = w35249 ^ w35240;
	assign w35201 = w35292 ^ w35293;
	assign w35248 = w35201 ^ w35202;
	assign w35247 = w35248 ^ w35230;
	assign w35289 = w35295 ^ w35247;
	assign w35291 = w35313 & w35304;
	assign w35286 = w35290 & w35289;
	assign w44846 = w35291 ^ w35297;
	assign w35241 = w44846 ^ w35226;
	assign w35287 = w35249 ^ w35241;
	assign w35203 = w35235 ^ w44846;
	assign w35246 = w940 ^ w35203;
	assign w35281 = w35286 ^ w35246;
	assign w44847 = w35291 ^ w35294;
	assign w35244 = w35292 ^ w44847;
	assign w35200 = w35295 ^ w35244;
	assign w35282 = w936 ^ w35200;
	assign w35280 = w35281 & w35282;
	assign w35278 = w35286 ^ w35280;
	assign w35199 = w35280 ^ w35244;
	assign w35198 = w35280 ^ w35297;
	assign w35193 = w35198 ^ w35294;
	assign w35204 = w35230 ^ w44847;
	assign w35288 = w35204 ^ w35229;
	assign w35279 = w35280 ^ w35288;
	assign w35285 = w35286 ^ w35288;
	assign w35284 = w35287 & w35285;
	assign w35283 = w35284 ^ w35246;
	assign w35195 = w35284 ^ w35296;
	assign w35191 = w35195 ^ w35231;
	assign w35194 = w942 ^ w35191;
	assign w35271 = w35193 ^ w35194;
	assign w35192 = w35284 ^ w35240;
	assign w35190 = w940 ^ w35191;
	assign w35277 = w35288 & w35278;
	assign w35275 = w35277 ^ w35285;
	assign w35274 = w35283 & w35275;
	assign w35239 = w35274 ^ w35249;
	assign w35273 = w35239 ^ w35241;
	assign w35197 = w35274 ^ w35298;
	assign w35270 = w35239 ^ w35192;
	assign w35265 = w35279 & w935;
	assign w35264 = w35270 & w35300;
	assign w35263 = w35273 & w35312;
	assign w35262 = w35283 & w35302;
	assign w35206 = w35262 ^ w35263;
	assign w35261 = w35271 & w35303;
	assign w35256 = w35279 & w35311;
	assign w35255 = w35270 & w35315;
	assign w35222 = w35264 ^ w35255;
	assign w35254 = w35273 & w35308;
	assign w35224 = w35262 ^ w35254;
	assign w35253 = w35283 & w35309;
	assign w35252 = w35271 & w35314;
	assign w44848 = w35263 ^ w35264;
	assign w44850 = w35277 ^ w35295;
	assign w35236 = w936 ^ w44850;
	assign w35189 = w35236 ^ w35197;
	assign w35196 = w35226 ^ w35189;
	assign w35272 = w35193 ^ w35196;
	assign w35259 = w35272 & w35304;
	assign w35237 = w35255 ^ w35259;
	assign w35215 = ~w35237;
	assign w35268 = w35189 ^ w35190;
	assign w35260 = w35268 & w35301;
	assign w35217 = w35260 ^ w35261;
	assign w35221 = w35260 ^ w35263;
	assign w35218 = ~w35221;
	assign w35214 = w35215 ^ w35253;
	assign w35251 = w35268 & w35316;
	assign w35250 = w35272 & w35313;
	assign w35216 = w35261 ^ w35250;
	assign w35212 = ~w35216;
	assign w43597 = w35251 ^ w35252;
	assign w35220 = w35224 ^ w43597;
	assign w35219 = w35215 ^ w35220;
	assign w35319 = w35218 ^ w35219;
	assign w48102 = ~w35319;
	assign w976 = w1741 ^ w48102;
	assign w1007 = w1772 ^ w976;
	assign w1039 = w1804 ^ w1007;
	assign w1071 = w1836 ^ w1039;
	assign w35276 = w35236 ^ w35199;
	assign w35266 = w35276 & w35305;
	assign w35257 = w35276 & w35307;
	assign w35233 = w35257 ^ w43597;
	assign w35245 = w35260 ^ w44848;
	assign w35211 = w35256 ^ w35245;
	assign w35208 = ~w35211;
	assign w35205 = w35261 ^ w35245;
	assign w35269 = w44850 ^ w35247;
	assign w35267 = w35269 & w35306;
	assign w35258 = w35269 & w35310;
	assign w35234 = w35258 ^ w35233;
	assign w35238 = w35266 ^ w35234;
	assign w35243 = w35267 ^ w35238;
	assign w48105 = w44848 ^ w35243;
	assign w979 = w1744 ^ w48105;
	assign w1010 = w1775 ^ w979;
	assign w1042 = w1807 ^ w1010;
	assign w1074 = w1839 ^ w1042;
	assign w35318 = w35243 ^ w35217;
	assign w35207 = w35265 ^ w35238;
	assign w48104 = w35206 ^ w35207;
	assign w978 = w1743 ^ w48104;
	assign w1009 = w1774 ^ w978;
	assign w1041 = w1806 ^ w1009;
	assign w1073 = w1838 ^ w1041;
	assign w35091 = w1071 ^ w1073;
	assign w48108 = w35234 ^ w35205;
	assign w982 = w1747 ^ w48108;
	assign w1013 = w1778 ^ w982;
	assign w1045 = w1810 ^ w1013;
	assign w1077 = w1842 ^ w1045;
	assign w35180 = w1074 ^ w1077;
	assign w35172 = w35091 ^ w35180;
	assign w35181 = w1077 ^ w1071;
	assign w48107 = ~w35318;
	assign w981 = w1746 ^ w48107;
	assign w1012 = w1777 ^ w981;
	assign w1044 = w1809 ^ w1012;
	assign w1076 = w1841 ^ w1044;
	assign w35094 = w1074 ^ w1076;
	assign w44849 = w35265 ^ w35267;
	assign w35223 = w44849 ^ w35220;
	assign w35320 = w35222 ^ w35223;
	assign w48101 = ~w35320;
	assign w975 = w1740 ^ w48101;
	assign w1006 = w1771 ^ w975;
	assign w1038 = w1803 ^ w1006;
	assign w1070 = w1835 ^ w1038;
	assign w35171 = w1070 ^ w35172;
	assign w35098 = w1070 ^ w1076;
	assign w35210 = w35214 ^ w44849;
	assign w35213 = w35252 ^ w35210;
	assign w35317 = w35212 ^ w35213;
	assign w35209 = w35233 ^ w35210;
	assign w48103 = w35208 ^ w35209;
	assign w977 = w1742 ^ w48103;
	assign w1008 = w1773 ^ w977;
	assign w1040 = w1805 ^ w1008;
	assign w1072 = w1837 ^ w1040;
	assign w35093 = w1072 ^ w35091;
	assign w35169 = w1076 ^ w35093;
	assign w35168 = w35098 ^ w35093;
	assign w35108 = w1071 ^ w1072;
	assign w35176 = w35180 ^ w35108;
	assign w35182 = w1072 ^ w1074;
	assign w35068 = w1073 ^ w1072;
	assign w35179 = w1077 ^ w1072;
	assign w35165 = w35172 & w35176;
	assign w35097 = w35165 ^ w35094;
	assign w35159 = w35180 & w35169;
	assign w35095 = w35159 ^ w35093;
	assign w35101 = w35097 ^ w35095;
	assign w35106 = w1077 ^ w35101;
	assign w48106 = ~w35317;
	assign w980 = w1745 ^ w48106;
	assign w1011 = w1776 ^ w980;
	assign w1043 = w1808 ^ w1011;
	assign w1075 = w1840 ^ w1043;
	assign w35166 = w1075 ^ w35093;
	assign w35092 = w1075 ^ w1077;
	assign w35167 = w35092 ^ w35182;
	assign w35175 = w35092 ^ w35098;
	assign w35173 = w35108 ^ w35175;
	assign w35178 = w1075 ^ w35098;
	assign w35174 = w1071 ^ w35178;
	assign w35054 = w35094 ^ w35092;
	assign w35170 = w35091 ^ w35054;
	assign w35053 = w35094 ^ w1075;
	assign w35177 = w1070 ^ w35053;
	assign w35164 = w35173 & w35171;
	assign w35163 = w35177 & w1070;
	assign w35162 = w35181 & w35166;
	assign w35096 = w35162 ^ w35092;
	assign w35161 = w35178 & w35174;
	assign w35160 = w35175 & w35168;
	assign w35158 = w35182 & w35167;
	assign w35115 = w35158 ^ w35164;
	assign w35156 = w35115 ^ w35106;
	assign w35067 = w35158 ^ w35159;
	assign w35114 = w35067 ^ w35068;
	assign w35113 = w35114 ^ w35096;
	assign w35155 = w35161 ^ w35113;
	assign w35157 = w35179 & w35170;
	assign w35152 = w35156 & w35155;
	assign w44840 = w35157 ^ w35160;
	assign w35070 = w35096 ^ w44840;
	assign w35154 = w35070 ^ w35095;
	assign w35151 = w35152 ^ w35154;
	assign w35110 = w35158 ^ w44840;
	assign w35066 = w35161 ^ w35110;
	assign w35148 = w1071 ^ w35066;
	assign w44843 = w35157 ^ w35163;
	assign w35069 = w35101 ^ w44843;
	assign w35112 = w1075 ^ w35069;
	assign w35147 = w35152 ^ w35112;
	assign w35146 = w35147 & w35148;
	assign w35145 = w35146 ^ w35154;
	assign w35144 = w35152 ^ w35146;
	assign w35065 = w35146 ^ w35110;
	assign w35064 = w35146 ^ w35163;
	assign w35059 = w35064 ^ w35160;
	assign w35143 = w35154 & w35144;
	assign w35141 = w35143 ^ w35151;
	assign w35131 = w35145 & w1070;
	assign w35122 = w35145 & w35177;
	assign w44842 = w35143 ^ w35161;
	assign w35135 = w44842 ^ w35113;
	assign w35133 = w35135 & w35172;
	assign w35124 = w35135 & w35176;
	assign w35102 = w1071 ^ w44842;
	assign w35142 = w35102 ^ w35065;
	assign w35132 = w35142 & w35171;
	assign w35123 = w35142 & w35173;
	assign w35107 = w44843 ^ w35092;
	assign w35153 = w35115 ^ w35107;
	assign w35150 = w35153 & w35151;
	assign w35149 = w35150 ^ w35112;
	assign w35061 = w35150 ^ w35162;
	assign w35057 = w35061 ^ w35097;
	assign w35060 = w1077 ^ w35057;
	assign w35137 = w35059 ^ w35060;
	assign w35058 = w35150 ^ w35106;
	assign w35056 = w1075 ^ w35057;
	assign w35140 = w35149 & w35141;
	assign w35105 = w35140 ^ w35115;
	assign w35139 = w35105 ^ w35107;
	assign w35063 = w35140 ^ w35164;
	assign w35055 = w35102 ^ w35063;
	assign w35062 = w35092 ^ w35055;
	assign w35138 = w35059 ^ w35062;
	assign w35136 = w35105 ^ w35058;
	assign w35134 = w35055 ^ w35056;
	assign w35130 = w35136 & w35166;
	assign w35129 = w35139 & w35178;
	assign w35128 = w35149 & w35168;
	assign w35072 = w35128 ^ w35129;
	assign w35127 = w35137 & w35169;
	assign w35126 = w35134 & w35167;
	assign w35087 = w35126 ^ w35129;
	assign w35084 = ~w35087;
	assign w35083 = w35126 ^ w35127;
	assign w35125 = w35138 & w35170;
	assign w35121 = w35136 & w35181;
	assign w35103 = w35121 ^ w35125;
	assign w35088 = w35130 ^ w35121;
	assign w35081 = ~w35103;
	assign w35120 = w35139 & w35174;
	assign w35090 = w35128 ^ w35120;
	assign w35119 = w35149 & w35175;
	assign w35080 = w35081 ^ w35119;
	assign w35118 = w35137 & w35180;
	assign w35117 = w35134 & w35182;
	assign w35116 = w35138 & w35179;
	assign w35082 = w35127 ^ w35116;
	assign w35078 = ~w35082;
	assign w44841 = w35117 ^ w35118;
	assign w35099 = w35123 ^ w44841;
	assign w35100 = w35124 ^ w35099;
	assign w35104 = w35132 ^ w35100;
	assign w35109 = w35133 ^ w35104;
	assign w35184 = w35109 ^ w35083;
	assign w35073 = w35131 ^ w35104;
	assign w48136 = w35072 ^ w35073;
	assign w1105 = w1870 ^ w48136;
	assign w48139 = ~w35184;
	assign w1108 = w1873 ^ w48139;
	assign w1140 = w885 ^ w1108;
	assign w1137 = w882 ^ w1105;
	assign w1172 = w917 ^ w1140;
	assign w1169 = w914 ^ w1137;
	assign w1201 = w946 ^ w1169;
	assign w1204 = w949 ^ w1172;
	assign w35086 = w35090 ^ w44841;
	assign w35085 = w35081 ^ w35086;
	assign w35185 = w35084 ^ w35085;
	assign w48134 = ~w35185;
	assign w1103 = w1868 ^ w48134;
	assign w1135 = w880 ^ w1103;
	assign w1167 = w912 ^ w1135;
	assign w1199 = w944 ^ w1167;
	assign w37771 = w1199 ^ w1201;
	assign w44844 = w35129 ^ w35130;
	assign w48137 = w44844 ^ w35109;
	assign w1106 = w1871 ^ w48137;
	assign w1138 = w883 ^ w1106;
	assign w1170 = w915 ^ w1138;
	assign w1202 = w947 ^ w1170;
	assign w37774 = w1202 ^ w1204;
	assign w35111 = w35126 ^ w44844;
	assign w35077 = w35122 ^ w35111;
	assign w35074 = ~w35077;
	assign w35071 = w35127 ^ w35111;
	assign w48140 = w35100 ^ w35071;
	assign w1109 = w1874 ^ w48140;
	assign w1141 = w886 ^ w1109;
	assign w1173 = w918 ^ w1141;
	assign w1205 = w950 ^ w1173;
	assign w37860 = w1202 ^ w1205;
	assign w37852 = w37771 ^ w37860;
	assign w37861 = w1205 ^ w1199;
	assign w44845 = w35131 ^ w35133;
	assign w35089 = w44845 ^ w35086;
	assign w35186 = w35088 ^ w35089;
	assign w48133 = ~w35186;
	assign w1102 = w1867 ^ w48133;
	assign w1134 = w879 ^ w1102;
	assign w1166 = w911 ^ w1134;
	assign w1198 = w943 ^ w1166;
	assign w37851 = w1198 ^ w37852;
	assign w37778 = w1198 ^ w1204;
	assign w35076 = w35080 ^ w44845;
	assign w35079 = w35118 ^ w35076;
	assign w35183 = w35078 ^ w35079;
	assign w35075 = w35099 ^ w35076;
	assign w48135 = w35074 ^ w35075;
	assign w1104 = w1869 ^ w48135;
	assign w48138 = ~w35183;
	assign w1107 = w1872 ^ w48138;
	assign w1139 = w884 ^ w1107;
	assign w1136 = w881 ^ w1104;
	assign w1171 = w916 ^ w1139;
	assign w1203 = w948 ^ w1171;
	assign w37772 = w1203 ^ w1205;
	assign w37855 = w37772 ^ w37778;
	assign w37858 = w1203 ^ w37778;
	assign w37854 = w1199 ^ w37858;
	assign w37734 = w37774 ^ w37772;
	assign w37850 = w37771 ^ w37734;
	assign w37733 = w37774 ^ w1203;
	assign w37857 = w1198 ^ w37733;
	assign w37843 = w37857 & w1198;
	assign w37841 = w37858 & w37854;
	assign w1168 = w913 ^ w1136;
	assign w1200 = w945 ^ w1168;
	assign w37773 = w1200 ^ w37771;
	assign w37849 = w1204 ^ w37773;
	assign w37846 = w1203 ^ w37773;
	assign w37848 = w37778 ^ w37773;
	assign w37788 = w1199 ^ w1200;
	assign w37853 = w37788 ^ w37855;
	assign w37856 = w37860 ^ w37788;
	assign w37862 = w1200 ^ w1202;
	assign w37847 = w37772 ^ w37862;
	assign w37748 = w1201 ^ w1200;
	assign w37859 = w1205 ^ w1200;
	assign w37845 = w37852 & w37856;
	assign w37777 = w37845 ^ w37774;
	assign w37844 = w37853 & w37851;
	assign w37842 = w37861 & w37846;
	assign w37776 = w37842 ^ w37772;
	assign w37840 = w37855 & w37848;
	assign w37839 = w37860 & w37849;
	assign w37775 = w37839 ^ w37773;
	assign w37781 = w37777 ^ w37775;
	assign w37786 = w1205 ^ w37781;
	assign w37838 = w37862 & w37847;
	assign w37795 = w37838 ^ w37844;
	assign w37836 = w37795 ^ w37786;
	assign w37747 = w37838 ^ w37839;
	assign w37794 = w37747 ^ w37748;
	assign w37793 = w37794 ^ w37776;
	assign w37835 = w37841 ^ w37793;
	assign w37837 = w37859 & w37850;
	assign w37832 = w37836 & w37835;
	assign w44953 = w37837 ^ w37843;
	assign w37749 = w37781 ^ w44953;
	assign w37792 = w1203 ^ w37749;
	assign w37827 = w37832 ^ w37792;
	assign w37787 = w44953 ^ w37772;
	assign w37833 = w37795 ^ w37787;
	assign w44954 = w37837 ^ w37840;
	assign w37790 = w37838 ^ w44954;
	assign w37746 = w37841 ^ w37790;
	assign w37828 = w1199 ^ w37746;
	assign w37826 = w37827 & w37828;
	assign w37824 = w37832 ^ w37826;
	assign w37745 = w37826 ^ w37790;
	assign w37744 = w37826 ^ w37843;
	assign w37739 = w37744 ^ w37840;
	assign w37750 = w37776 ^ w44954;
	assign w37834 = w37750 ^ w37775;
	assign w37825 = w37826 ^ w37834;
	assign w37831 = w37832 ^ w37834;
	assign w37830 = w37833 & w37831;
	assign w37829 = w37830 ^ w37792;
	assign w37741 = w37830 ^ w37842;
	assign w37737 = w37741 ^ w37777;
	assign w37740 = w1205 ^ w37737;
	assign w37817 = w37739 ^ w37740;
	assign w37738 = w37830 ^ w37786;
	assign w37736 = w1203 ^ w37737;
	assign w37823 = w37834 & w37824;
	assign w37821 = w37823 ^ w37831;
	assign w37820 = w37829 & w37821;
	assign w37785 = w37820 ^ w37795;
	assign w37819 = w37785 ^ w37787;
	assign w37743 = w37820 ^ w37844;
	assign w37816 = w37785 ^ w37738;
	assign w37811 = w37825 & w1198;
	assign w37810 = w37816 & w37846;
	assign w37809 = w37819 & w37858;
	assign w37808 = w37829 & w37848;
	assign w37752 = w37808 ^ w37809;
	assign w37807 = w37817 & w37849;
	assign w37802 = w37825 & w37857;
	assign w37801 = w37816 & w37861;
	assign w37768 = w37810 ^ w37801;
	assign w37800 = w37819 & w37854;
	assign w37770 = w37808 ^ w37800;
	assign w37799 = w37829 & w37855;
	assign w37798 = w37817 & w37860;
	assign w44956 = w37809 ^ w37810;
	assign w44958 = w37823 ^ w37841;
	assign w37815 = w44958 ^ w37793;
	assign w37804 = w37815 & w37856;
	assign w37813 = w37815 & w37852;
	assign w44957 = w37811 ^ w37813;
	assign w37782 = w1199 ^ w44958;
	assign w37822 = w37782 ^ w37745;
	assign w37735 = w37782 ^ w37743;
	assign w37742 = w37772 ^ w37735;
	assign w37818 = w37739 ^ w37742;
	assign w37814 = w37735 ^ w37736;
	assign w37812 = w37822 & w37851;
	assign w37806 = w37814 & w37847;
	assign w37791 = w37806 ^ w44956;
	assign w37767 = w37806 ^ w37809;
	assign w37764 = ~w37767;
	assign w37763 = w37806 ^ w37807;
	assign w37757 = w37802 ^ w37791;
	assign w37754 = ~w37757;
	assign w37751 = w37807 ^ w37791;
	assign w37805 = w37818 & w37850;
	assign w37783 = w37801 ^ w37805;
	assign w37761 = ~w37783;
	assign w37760 = w37761 ^ w37799;
	assign w37756 = w37760 ^ w44957;
	assign w37759 = w37798 ^ w37756;
	assign w37803 = w37822 & w37853;
	assign w37797 = w37814 & w37862;
	assign w37796 = w37818 & w37859;
	assign w37762 = w37807 ^ w37796;
	assign w37758 = ~w37762;
	assign w37863 = w37758 ^ w37759;
	assign w48178 = ~w37863;
	assign w1242 = w987 ^ w48178;
	assign w1274 = w1019 ^ w1242;
	assign w1306 = w1051 ^ w1274;
	assign w1338 = w1083 ^ w1306;
	assign w44955 = w37797 ^ w37798;
	assign w37779 = w37803 ^ w44955;
	assign w37755 = w37779 ^ w37756;
	assign w48175 = w37754 ^ w37755;
	assign w37780 = w37804 ^ w37779;
	assign w48180 = w37780 ^ w37751;
	assign w37784 = w37812 ^ w37780;
	assign w37753 = w37811 ^ w37784;
	assign w48176 = w37752 ^ w37753;
	assign w37789 = w37813 ^ w37784;
	assign w37864 = w37789 ^ w37763;
	assign w48179 = ~w37864;
	assign w1243 = w988 ^ w48179;
	assign w1275 = w1020 ^ w1243;
	assign w1307 = w1052 ^ w1275;
	assign w1339 = w1084 ^ w1307;
	assign w1244 = w989 ^ w48180;
	assign w1276 = w1021 ^ w1244;
	assign w1308 = w1053 ^ w1276;
	assign w1340 = w1085 ^ w1308;
	assign w37638 = w1338 ^ w1340;
	assign w48177 = w44956 ^ w37789;
	assign w2046 = w986 ^ w48177;
	assign w37766 = w37770 ^ w44955;
	assign w37769 = w44957 ^ w37766;
	assign w37866 = w37768 ^ w37769;
	assign w37765 = w37761 ^ w37766;
	assign w37865 = w37764 ^ w37765;
	assign w48173 = ~w37866;
	assign w1238 = w983 ^ w48173;
	assign w1269 = w1014 ^ w1238;
	assign w1301 = w1046 ^ w1269;
	assign w1333 = w1078 ^ w1301;
	assign w37644 = w1333 ^ w1339;
	assign w37721 = w37638 ^ w37644;
	assign w37724 = w1338 ^ w37644;
	assign w48174 = ~w37865;
	assign w1239 = w984 ^ w48174;
	assign w1270 = w1015 ^ w1239;
	assign w1302 = w1047 ^ w1270;
	assign w1334 = w1079 ^ w1302;
	assign w37720 = w1334 ^ w37724;
	assign w37727 = w1340 ^ w1334;
	assign w37707 = w37724 & w37720;
	assign w44982 = w38507 ^ w38513;
	assign w38457 = w44982 ^ w38442;
	assign w38503 = w38465 ^ w38457;
	assign w38419 = w38451 ^ w44982;
	assign w38462 = w1593 ^ w38419;
	assign w38497 = w38502 ^ w38462;
	assign w44983 = w38507 ^ w38510;
	assign w38460 = w38508 ^ w44983;
	assign w38416 = w38511 ^ w38460;
	assign w38498 = w1589 ^ w38416;
	assign w38496 = w38497 & w38498;
	assign w38415 = w38496 ^ w38460;
	assign w38414 = w38496 ^ w38513;
	assign w38409 = w38414 ^ w38510;
	assign w38494 = w38502 ^ w38496;
	assign w38420 = w38446 ^ w44983;
	assign w38504 = w38420 ^ w38445;
	assign w38495 = w38496 ^ w38504;
	assign w38501 = w38502 ^ w38504;
	assign w38500 = w38503 & w38501;
	assign w38499 = w38500 ^ w38462;
	assign w38411 = w38500 ^ w38512;
	assign w38407 = w38411 ^ w38447;
	assign w38410 = w1595 ^ w38407;
	assign w38487 = w38409 ^ w38410;
	assign w38408 = w38500 ^ w38456;
	assign w38406 = w1593 ^ w38407;
	assign w38493 = w38504 & w38494;
	assign w38491 = w38493 ^ w38501;
	assign w38490 = w38499 & w38491;
	assign w38455 = w38490 ^ w38465;
	assign w38489 = w38455 ^ w38457;
	assign w38413 = w38490 ^ w38514;
	assign w38486 = w38455 ^ w38408;
	assign w38481 = w38495 & w1588;
	assign w38480 = w38486 & w38516;
	assign w38479 = w38489 & w38528;
	assign w38478 = w38499 & w38518;
	assign w38422 = w38478 ^ w38479;
	assign w38477 = w38487 & w38519;
	assign w38472 = w38495 & w38527;
	assign w38471 = w38486 & w38531;
	assign w38438 = w38480 ^ w38471;
	assign w38470 = w38489 & w38524;
	assign w38440 = w38478 ^ w38470;
	assign w38469 = w38499 & w38525;
	assign w38468 = w38487 & w38530;
	assign w44984 = w38479 ^ w38480;
	assign w44986 = w38493 ^ w38511;
	assign w38452 = w1589 ^ w44986;
	assign w38492 = w38452 ^ w38415;
	assign w38473 = w38492 & w38523;
	assign w38482 = w38492 & w38521;
	assign w38405 = w38452 ^ w38413;
	assign w38412 = w38442 ^ w38405;
	assign w38488 = w38409 ^ w38412;
	assign w38475 = w38488 & w38520;
	assign w38453 = w38471 ^ w38475;
	assign w38431 = ~w38453;
	assign w38430 = w38431 ^ w38469;
	assign w38484 = w38405 ^ w38406;
	assign w38467 = w38484 & w38532;
	assign w38466 = w38488 & w38529;
	assign w38432 = w38477 ^ w38466;
	assign w38428 = ~w38432;
	assign w43605 = w38467 ^ w38468;
	assign w38449 = w38473 ^ w43605;
	assign w38436 = w38440 ^ w43605;
	assign w38435 = w38431 ^ w38436;
	assign w38476 = w38484 & w38517;
	assign w38437 = w38476 ^ w38479;
	assign w38434 = ~w38437;
	assign w38535 = w38434 ^ w38435;
	assign w48014 = ~w38535;
	assign w1621 = w2035 ^ w48014;
	assign w1653 = w1398 ^ w1621;
	assign w1685 = w1430 ^ w1653;
	assign w1717 = w1462 ^ w1685;
	assign w38433 = w38476 ^ w38477;
	assign w38461 = w38476 ^ w44984;
	assign w38427 = w38472 ^ w38461;
	assign w38424 = ~w38427;
	assign w38421 = w38477 ^ w38461;
	assign w38485 = w44986 ^ w38463;
	assign w38483 = w38485 & w38522;
	assign w38474 = w38485 & w38526;
	assign w38450 = w38474 ^ w38449;
	assign w38454 = w38482 ^ w38450;
	assign w38459 = w38483 ^ w38454;
	assign w48017 = w44984 ^ w38459;
	assign w1624 = w2038 ^ w48017;
	assign w1656 = w1401 ^ w1624;
	assign w1688 = w1433 ^ w1656;
	assign w1720 = w1465 ^ w1688;
	assign w38534 = w38459 ^ w38433;
	assign w38423 = w38481 ^ w38454;
	assign w48016 = w38422 ^ w38423;
	assign w1623 = w2037 ^ w48016;
	assign w1655 = w1400 ^ w1623;
	assign w1687 = w1432 ^ w1655;
	assign w1719 = w1464 ^ w1687;
	assign w37101 = w1717 ^ w1719;
	assign w48020 = w38450 ^ w38421;
	assign w1627 = w2041 ^ w48020;
	assign w1659 = w1404 ^ w1627;
	assign w1691 = w1436 ^ w1659;
	assign w1723 = w1468 ^ w1691;
	assign w37190 = w1720 ^ w1723;
	assign w37182 = w37101 ^ w37190;
	assign w37191 = w1723 ^ w1717;
	assign w48019 = ~w38534;
	assign w1626 = w2040 ^ w48019;
	assign w1658 = w1403 ^ w1626;
	assign w1690 = w1435 ^ w1658;
	assign w1722 = w1467 ^ w1690;
	assign w37104 = w1720 ^ w1722;
	assign w44985 = w38481 ^ w38483;
	assign w38439 = w44985 ^ w38436;
	assign w38536 = w38438 ^ w38439;
	assign w48013 = ~w38536;
	assign w1620 = w2034 ^ w48013;
	assign w1652 = w1397 ^ w1620;
	assign w1684 = w1429 ^ w1652;
	assign w1716 = w1461 ^ w1684;
	assign w37108 = w1716 ^ w1722;
	assign w37181 = w1716 ^ w37182;
	assign w38426 = w38430 ^ w44985;
	assign w38429 = w38468 ^ w38426;
	assign w38533 = w38428 ^ w38429;
	assign w38425 = w38449 ^ w38426;
	assign w48015 = w38424 ^ w38425;
	assign w1622 = w2036 ^ w48015;
	assign w1654 = w1399 ^ w1622;
	assign w1686 = w1431 ^ w1654;
	assign w1718 = w1463 ^ w1686;
	assign w37103 = w1718 ^ w37101;
	assign w37179 = w1722 ^ w37103;
	assign w37178 = w37108 ^ w37103;
	assign w37118 = w1717 ^ w1718;
	assign w37186 = w37190 ^ w37118;
	assign w37192 = w1718 ^ w1720;
	assign w37078 = w1719 ^ w1718;
	assign w37189 = w1723 ^ w1718;
	assign w37175 = w37182 & w37186;
	assign w37107 = w37175 ^ w37104;
	assign w37169 = w37190 & w37179;
	assign w37105 = w37169 ^ w37103;
	assign w37111 = w37107 ^ w37105;
	assign w37116 = w1723 ^ w37111;
	assign w48018 = ~w38533;
	assign w1625 = w2039 ^ w48018;
	assign w1657 = w1402 ^ w1625;
	assign w1689 = w1434 ^ w1657;
	assign w1721 = w1466 ^ w1689;
	assign w37176 = w1721 ^ w37103;
	assign w37102 = w1721 ^ w1723;
	assign w37177 = w37102 ^ w37192;
	assign w37185 = w37102 ^ w37108;
	assign w37183 = w37118 ^ w37185;
	assign w37188 = w1721 ^ w37108;
	assign w37184 = w1717 ^ w37188;
	assign w37064 = w37104 ^ w37102;
	assign w37180 = w37101 ^ w37064;
	assign w37063 = w37104 ^ w1721;
	assign w37187 = w1716 ^ w37063;
	assign w37174 = w37183 & w37181;
	assign w37173 = w37187 & w1716;
	assign w37172 = w37191 & w37176;
	assign w37106 = w37172 ^ w37102;
	assign w37171 = w37188 & w37184;
	assign w37170 = w37185 & w37178;
	assign w37168 = w37192 & w37177;
	assign w37125 = w37168 ^ w37174;
	assign w37166 = w37125 ^ w37116;
	assign w37077 = w37168 ^ w37169;
	assign w37124 = w37077 ^ w37078;
	assign w37123 = w37124 ^ w37106;
	assign w37165 = w37171 ^ w37123;
	assign w37167 = w37189 & w37180;
	assign w37162 = w37166 & w37165;
	assign w44925 = w37167 ^ w37170;
	assign w37080 = w37106 ^ w44925;
	assign w37164 = w37080 ^ w37105;
	assign w37161 = w37162 ^ w37164;
	assign w37120 = w37168 ^ w44925;
	assign w37076 = w37171 ^ w37120;
	assign w37158 = w1717 ^ w37076;
	assign w44928 = w37167 ^ w37173;
	assign w37079 = w37111 ^ w44928;
	assign w37122 = w1721 ^ w37079;
	assign w37157 = w37162 ^ w37122;
	assign w37156 = w37157 & w37158;
	assign w37154 = w37162 ^ w37156;
	assign w37075 = w37156 ^ w37120;
	assign w37074 = w37156 ^ w37173;
	assign w37069 = w37074 ^ w37170;
	assign w37153 = w37164 & w37154;
	assign w37151 = w37153 ^ w37161;
	assign w44927 = w37153 ^ w37171;
	assign w37145 = w44927 ^ w37123;
	assign w37134 = w37145 & w37186;
	assign w37143 = w37145 & w37182;
	assign w37112 = w1717 ^ w44927;
	assign w37152 = w37112 ^ w37075;
	assign w37142 = w37152 & w37181;
	assign w37133 = w37152 & w37183;
	assign w37155 = w37156 ^ w37164;
	assign w37141 = w37155 & w1716;
	assign w37132 = w37155 & w37187;
	assign w37117 = w44928 ^ w37102;
	assign w37163 = w37125 ^ w37117;
	assign w37160 = w37163 & w37161;
	assign w37159 = w37160 ^ w37122;
	assign w37071 = w37160 ^ w37172;
	assign w37067 = w37071 ^ w37107;
	assign w37070 = w1723 ^ w37067;
	assign w37147 = w37069 ^ w37070;
	assign w37068 = w37160 ^ w37116;
	assign w37066 = w1721 ^ w37067;
	assign w37150 = w37159 & w37151;
	assign w37115 = w37150 ^ w37125;
	assign w37149 = w37115 ^ w37117;
	assign w37073 = w37150 ^ w37174;
	assign w37065 = w37112 ^ w37073;
	assign w37072 = w37102 ^ w37065;
	assign w37148 = w37069 ^ w37072;
	assign w37146 = w37115 ^ w37068;
	assign w37144 = w37065 ^ w37066;
	assign w37140 = w37146 & w37176;
	assign w37139 = w37149 & w37188;
	assign w37138 = w37159 & w37178;
	assign w37082 = w37138 ^ w37139;
	assign w37137 = w37147 & w37179;
	assign w37136 = w37144 & w37177;
	assign w37097 = w37136 ^ w37139;
	assign w37094 = ~w37097;
	assign w37093 = w37136 ^ w37137;
	assign w37135 = w37148 & w37180;
	assign w37131 = w37146 & w37191;
	assign w37113 = w37131 ^ w37135;
	assign w37098 = w37140 ^ w37131;
	assign w37091 = ~w37113;
	assign w37130 = w37149 & w37184;
	assign w37100 = w37138 ^ w37130;
	assign w37129 = w37159 & w37185;
	assign w37090 = w37091 ^ w37129;
	assign w37128 = w37147 & w37190;
	assign w37127 = w37144 & w37192;
	assign w37126 = w37148 & w37189;
	assign w37092 = w37137 ^ w37126;
	assign w37088 = ~w37092;
	assign w44926 = w37127 ^ w37128;
	assign w37096 = w37100 ^ w44926;
	assign w37095 = w37091 ^ w37096;
	assign w37195 = w37094 ^ w37095;
	assign w48022 = ~w37195;
	assign w1725 = w1470 ^ w48022;
	assign w1756 = w1501 ^ w1725;
	assign w1788 = w1533 ^ w1756;
	assign w1820 = w1565 ^ w1788;
	assign w37109 = w37133 ^ w44926;
	assign w37110 = w37134 ^ w37109;
	assign w37114 = w37142 ^ w37110;
	assign w37119 = w37143 ^ w37114;
	assign w37194 = w37119 ^ w37093;
	assign w37083 = w37141 ^ w37114;
	assign w48024 = w37082 ^ w37083;
	assign w1727 = w1472 ^ w48024;
	assign w1758 = w1503 ^ w1727;
	assign w1790 = w1535 ^ w1758;
	assign w1822 = w1567 ^ w1790;
	assign w36967 = w1820 ^ w1822;
	assign w48027 = ~w37194;
	assign w1730 = w1475 ^ w48027;
	assign w1761 = w1506 ^ w1730;
	assign w1793 = w1538 ^ w1761;
	assign w1825 = w1570 ^ w1793;
	assign w44929 = w37139 ^ w37140;
	assign w48025 = w44929 ^ w37119;
	assign w1728 = w1473 ^ w48025;
	assign w1759 = w1504 ^ w1728;
	assign w1791 = w1536 ^ w1759;
	assign w1823 = w1568 ^ w1791;
	assign w36970 = w1823 ^ w1825;
	assign w37121 = w37136 ^ w44929;
	assign w37087 = w37132 ^ w37121;
	assign w37084 = ~w37087;
	assign w37081 = w37137 ^ w37121;
	assign w48028 = w37110 ^ w37081;
	assign w1731 = w1476 ^ w48028;
	assign w1762 = w1507 ^ w1731;
	assign w1794 = w1539 ^ w1762;
	assign w1826 = w1571 ^ w1794;
	assign w37056 = w1823 ^ w1826;
	assign w37048 = w36967 ^ w37056;
	assign w37057 = w1826 ^ w1820;
	assign w44930 = w37141 ^ w37143;
	assign w37099 = w44930 ^ w37096;
	assign w37196 = w37098 ^ w37099;
	assign w48021 = ~w37196;
	assign w1724 = w1469 ^ w48021;
	assign w1755 = w1500 ^ w1724;
	assign w1787 = w1532 ^ w1755;
	assign w1819 = w1564 ^ w1787;
	assign w37047 = w1819 ^ w37048;
	assign w36974 = w1819 ^ w1825;
	assign w37086 = w37090 ^ w44930;
	assign w37089 = w37128 ^ w37086;
	assign w37193 = w37088 ^ w37089;
	assign w37085 = w37109 ^ w37086;
	assign w48023 = w37084 ^ w37085;
	assign w1726 = w1471 ^ w48023;
	assign w1757 = w1502 ^ w1726;
	assign w1789 = w1534 ^ w1757;
	assign w1821 = w1566 ^ w1789;
	assign w36969 = w1821 ^ w36967;
	assign w37045 = w1825 ^ w36969;
	assign w37044 = w36974 ^ w36969;
	assign w36984 = w1820 ^ w1821;
	assign w37052 = w37056 ^ w36984;
	assign w37058 = w1821 ^ w1823;
	assign w36944 = w1822 ^ w1821;
	assign w37055 = w1826 ^ w1821;
	assign w37041 = w37048 & w37052;
	assign w36973 = w37041 ^ w36970;
	assign w37035 = w37056 & w37045;
	assign w36971 = w37035 ^ w36969;
	assign w36977 = w36973 ^ w36971;
	assign w36982 = w1826 ^ w36977;
	assign w48026 = ~w37193;
	assign w1729 = w1474 ^ w48026;
	assign w1760 = w1505 ^ w1729;
	assign w1792 = w1537 ^ w1760;
	assign w1824 = w1569 ^ w1792;
	assign w37042 = w1824 ^ w36969;
	assign w36968 = w1824 ^ w1826;
	assign w37043 = w36968 ^ w37058;
	assign w37051 = w36968 ^ w36974;
	assign w37049 = w36984 ^ w37051;
	assign w37054 = w1824 ^ w36974;
	assign w37050 = w1820 ^ w37054;
	assign w36930 = w36970 ^ w36968;
	assign w37046 = w36967 ^ w36930;
	assign w36929 = w36970 ^ w1824;
	assign w37053 = w1819 ^ w36929;
	assign w37040 = w37049 & w37047;
	assign w37039 = w37053 & w1819;
	assign w37038 = w37057 & w37042;
	assign w36972 = w37038 ^ w36968;
	assign w37037 = w37054 & w37050;
	assign w37036 = w37051 & w37044;
	assign w37034 = w37058 & w37043;
	assign w36991 = w37034 ^ w37040;
	assign w37032 = w36991 ^ w36982;
	assign w36943 = w37034 ^ w37035;
	assign w36990 = w36943 ^ w36944;
	assign w36989 = w36990 ^ w36972;
	assign w37031 = w37037 ^ w36989;
	assign w37033 = w37055 & w37046;
	assign w37028 = w37032 & w37031;
	assign w44919 = w37033 ^ w37039;
	assign w36945 = w36977 ^ w44919;
	assign w36988 = w1824 ^ w36945;
	assign w37023 = w37028 ^ w36988;
	assign w36983 = w44919 ^ w36968;
	assign w37029 = w36991 ^ w36983;
	assign w44920 = w37033 ^ w37036;
	assign w36986 = w37034 ^ w44920;
	assign w36942 = w37037 ^ w36986;
	assign w37024 = w1820 ^ w36942;
	assign w37022 = w37023 & w37024;
	assign w36941 = w37022 ^ w36986;
	assign w37020 = w37028 ^ w37022;
	assign w36940 = w37022 ^ w37039;
	assign w36935 = w36940 ^ w37036;
	assign w36946 = w36972 ^ w44920;
	assign w37030 = w36946 ^ w36971;
	assign w37021 = w37022 ^ w37030;
	assign w37027 = w37028 ^ w37030;
	assign w37026 = w37029 & w37027;
	assign w37025 = w37026 ^ w36988;
	assign w36937 = w37026 ^ w37038;
	assign w36933 = w36937 ^ w36973;
	assign w36936 = w1826 ^ w36933;
	assign w37013 = w36935 ^ w36936;
	assign w36934 = w37026 ^ w36982;
	assign w36932 = w1824 ^ w36933;
	assign w37019 = w37030 & w37020;
	assign w37017 = w37019 ^ w37027;
	assign w37016 = w37025 & w37017;
	assign w36981 = w37016 ^ w36991;
	assign w37015 = w36981 ^ w36983;
	assign w36939 = w37016 ^ w37040;
	assign w37012 = w36981 ^ w36934;
	assign w37007 = w37021 & w1819;
	assign w37006 = w37012 & w37042;
	assign w37005 = w37015 & w37054;
	assign w37004 = w37025 & w37044;
	assign w36948 = w37004 ^ w37005;
	assign w37003 = w37013 & w37045;
	assign w36998 = w37021 & w37053;
	assign w36997 = w37012 & w37057;
	assign w36964 = w37006 ^ w36997;
	assign w36996 = w37015 & w37050;
	assign w36966 = w37004 ^ w36996;
	assign w36995 = w37025 & w37051;
	assign w36994 = w37013 & w37056;
	assign w44922 = w37005 ^ w37006;
	assign w44924 = w37019 ^ w37037;
	assign w37011 = w44924 ^ w36989;
	assign w37009 = w37011 & w37048;
	assign w44923 = w37007 ^ w37009;
	assign w37000 = w37011 & w37052;
	assign w36978 = w1820 ^ w44924;
	assign w37018 = w36978 ^ w36941;
	assign w36931 = w36978 ^ w36939;
	assign w36938 = w36968 ^ w36931;
	assign w37014 = w36935 ^ w36938;
	assign w37010 = w36931 ^ w36932;
	assign w37008 = w37018 & w37047;
	assign w37002 = w37010 & w37043;
	assign w36987 = w37002 ^ w44922;
	assign w36963 = w37002 ^ w37005;
	assign w36960 = ~w36963;
	assign w36959 = w37002 ^ w37003;
	assign w36953 = w36998 ^ w36987;
	assign w36950 = ~w36953;
	assign w36947 = w37003 ^ w36987;
	assign w37001 = w37014 & w37046;
	assign w36979 = w36997 ^ w37001;
	assign w36957 = ~w36979;
	assign w36956 = w36957 ^ w36995;
	assign w36952 = w36956 ^ w44923;
	assign w36955 = w36994 ^ w36952;
	assign w36999 = w37018 & w37049;
	assign w36993 = w37010 & w37058;
	assign w36992 = w37014 & w37055;
	assign w36958 = w37003 ^ w36992;
	assign w36954 = ~w36958;
	assign w37059 = w36954 ^ w36955;
	assign w48058 = ~w37059;
	assign w1856 = w1601 ^ w48058;
	assign w868 = w1633 ^ w1856;
	assign w900 = w1665 ^ w868;
	assign w932 = w1697 ^ w900;
	assign w44921 = w36993 ^ w36994;
	assign w36962 = w36966 ^ w44921;
	assign w36965 = w44923 ^ w36962;
	assign w37062 = w36964 ^ w36965;
	assign w36961 = w36957 ^ w36962;
	assign w37061 = w36960 ^ w36961;
	assign w48054 = ~w37061;
	assign w1852 = w1597 ^ w48054;
	assign w864 = w1629 ^ w1852;
	assign w896 = w1661 ^ w864;
	assign w928 = w1693 ^ w896;
	assign w48053 = ~w37062;
	assign w1851 = w1596 ^ w48053;
	assign w863 = w1628 ^ w1851;
	assign w895 = w1660 ^ w863;
	assign w927 = w1692 ^ w895;
	assign w36975 = w36999 ^ w44921;
	assign w36976 = w37000 ^ w36975;
	assign w36980 = w37008 ^ w36976;
	assign w36985 = w37009 ^ w36980;
	assign w48057 = w44922 ^ w36985;
	assign w1855 = w1600 ^ w48057;
	assign w867 = w1632 ^ w1855;
	assign w899 = w1664 ^ w867;
	assign w931 = w1696 ^ w899;
	assign w37060 = w36985 ^ w36959;
	assign w36951 = w36975 ^ w36952;
	assign w48055 = w36950 ^ w36951;
	assign w1853 = w1598 ^ w48055;
	assign w865 = w1630 ^ w1853;
	assign w897 = w1662 ^ w865;
	assign w929 = w1694 ^ w897;
	assign w22914 = w928 ^ w929;
	assign w22988 = w929 ^ w931;
	assign w36949 = w37007 ^ w36980;
	assign w48056 = w36948 ^ w36949;
	assign w1854 = w1599 ^ w48056;
	assign w866 = w1631 ^ w1854;
	assign w898 = w1663 ^ w866;
	assign w930 = w1695 ^ w898;
	assign w22897 = w928 ^ w930;
	assign w22899 = w929 ^ w22897;
	assign w22972 = w932 ^ w22899;
	assign w22874 = w930 ^ w929;
	assign w48060 = w36976 ^ w36947;
	assign w1858 = w1603 ^ w48060;
	assign w870 = w1635 ^ w1858;
	assign w902 = w1667 ^ w870;
	assign w934 = w1699 ^ w902;
	assign w22898 = w932 ^ w934;
	assign w22973 = w22898 ^ w22988;
	assign w22986 = w931 ^ w934;
	assign w22982 = w22986 ^ w22914;
	assign w22978 = w22897 ^ w22986;
	assign w22977 = w927 ^ w22978;
	assign w22987 = w934 ^ w928;
	assign w22985 = w934 ^ w929;
	assign w22971 = w22978 & w22982;
	assign w22968 = w22987 & w22972;
	assign w22902 = w22968 ^ w22898;
	assign w22964 = w22988 & w22973;
	assign w48059 = ~w37060;
	assign w1857 = w1602 ^ w48059;
	assign w869 = w1634 ^ w1857;
	assign w901 = w1666 ^ w869;
	assign w933 = w1698 ^ w901;
	assign w22975 = w933 ^ w22899;
	assign w22900 = w931 ^ w933;
	assign w22903 = w22971 ^ w22900;
	assign w22904 = w927 ^ w933;
	assign w22974 = w22904 ^ w22899;
	assign w22981 = w22898 ^ w22904;
	assign w22979 = w22914 ^ w22981;
	assign w22984 = w932 ^ w22904;
	assign w22980 = w928 ^ w22984;
	assign w22860 = w22900 ^ w22898;
	assign w22976 = w22897 ^ w22860;
	assign w22859 = w22900 ^ w932;
	assign w22983 = w927 ^ w22859;
	assign w22970 = w22979 & w22977;
	assign w22921 = w22964 ^ w22970;
	assign w22969 = w22983 & w927;
	assign w22967 = w22984 & w22980;
	assign w22966 = w22981 & w22974;
	assign w22965 = w22986 & w22975;
	assign w22901 = w22965 ^ w22899;
	assign w22907 = w22903 ^ w22901;
	assign w22912 = w934 ^ w22907;
	assign w22962 = w22921 ^ w22912;
	assign w22873 = w22964 ^ w22965;
	assign w22920 = w22873 ^ w22874;
	assign w22919 = w22920 ^ w22902;
	assign w22961 = w22967 ^ w22919;
	assign w22963 = w22985 & w22976;
	assign w22958 = w22962 & w22961;
	assign w44329 = w22963 ^ w22969;
	assign w22913 = w44329 ^ w22898;
	assign w22959 = w22921 ^ w22913;
	assign w22875 = w22907 ^ w44329;
	assign w22918 = w932 ^ w22875;
	assign w22953 = w22958 ^ w22918;
	assign w44330 = w22963 ^ w22966;
	assign w22916 = w22964 ^ w44330;
	assign w22872 = w22967 ^ w22916;
	assign w22954 = w928 ^ w22872;
	assign w22952 = w22953 & w22954;
	assign w22871 = w22952 ^ w22916;
	assign w22870 = w22952 ^ w22969;
	assign w22865 = w22870 ^ w22966;
	assign w22950 = w22958 ^ w22952;
	assign w22876 = w22902 ^ w44330;
	assign w22960 = w22876 ^ w22901;
	assign w22951 = w22952 ^ w22960;
	assign w22957 = w22958 ^ w22960;
	assign w22956 = w22959 & w22957;
	assign w22955 = w22956 ^ w22918;
	assign w22867 = w22956 ^ w22968;
	assign w22863 = w22867 ^ w22903;
	assign w22866 = w934 ^ w22863;
	assign w22943 = w22865 ^ w22866;
	assign w22864 = w22956 ^ w22912;
	assign w22862 = w932 ^ w22863;
	assign w22949 = w22960 & w22950;
	assign w22947 = w22949 ^ w22957;
	assign w22946 = w22955 & w22947;
	assign w22911 = w22946 ^ w22921;
	assign w22945 = w22911 ^ w22913;
	assign w22869 = w22946 ^ w22970;
	assign w22942 = w22911 ^ w22864;
	assign w22937 = w22951 & w927;
	assign w22936 = w22942 & w22972;
	assign w22935 = w22945 & w22984;
	assign w22934 = w22955 & w22974;
	assign w22878 = w22934 ^ w22935;
	assign w22933 = w22943 & w22975;
	assign w22928 = w22951 & w22983;
	assign w22927 = w22942 & w22987;
	assign w22894 = w22936 ^ w22927;
	assign w22926 = w22945 & w22980;
	assign w22896 = w22934 ^ w22926;
	assign w22925 = w22955 & w22981;
	assign w22924 = w22943 & w22986;
	assign w44331 = w22935 ^ w22936;
	assign w44333 = w22949 ^ w22967;
	assign w22908 = w928 ^ w44333;
	assign w22948 = w22908 ^ w22871;
	assign w22929 = w22948 & w22979;
	assign w22938 = w22948 & w22977;
	assign w22861 = w22908 ^ w22869;
	assign w22868 = w22898 ^ w22861;
	assign w22944 = w22865 ^ w22868;
	assign w22931 = w22944 & w22976;
	assign w22909 = w22927 ^ w22931;
	assign w22887 = ~w22909;
	assign w22886 = w22887 ^ w22925;
	assign w22940 = w22861 ^ w22862;
	assign w22923 = w22940 & w22988;
	assign w22922 = w22944 & w22985;
	assign w22888 = w22933 ^ w22922;
	assign w22884 = ~w22888;
	assign w43562 = w22923 ^ w22924;
	assign w22905 = w22929 ^ w43562;
	assign w22892 = w22896 ^ w43562;
	assign w22891 = w22887 ^ w22892;
	assign w22932 = w22940 & w22973;
	assign w22889 = w22932 ^ w22933;
	assign w22917 = w22932 ^ w44331;
	assign w22883 = w22928 ^ w22917;
	assign w22880 = ~w22883;
	assign w22877 = w22933 ^ w22917;
	assign w22893 = w22932 ^ w22935;
	assign w22890 = ~w22893;
	assign w22991 = w22890 ^ w22891;
	assign w48094 = ~w22991;
	assign w968 = w1733 ^ w48094;
	assign w999 = w1764 ^ w968;
	assign w1031 = w1796 ^ w999;
	assign w1063 = w1828 ^ w1031;
	assign w22941 = w44333 ^ w22919;
	assign w22939 = w22941 & w22978;
	assign w22930 = w22941 & w22982;
	assign w22906 = w22930 ^ w22905;
	assign w22910 = w22938 ^ w22906;
	assign w22915 = w22939 ^ w22910;
	assign w48097 = w44331 ^ w22915;
	assign w22990 = w22915 ^ w22889;
	assign w22879 = w22937 ^ w22910;
	assign w48096 = w22878 ^ w22879;
	assign w48100 = w22906 ^ w22877;
	assign w48099 = ~w22990;
	assign w970 = w1735 ^ w48096;
	assign w974 = w1739 ^ w48100;
	assign w971 = w1736 ^ w48097;
	assign w973 = w1738 ^ w48099;
	assign w1005 = w1770 ^ w974;
	assign w1037 = w1802 ^ w1005;
	assign w1004 = w1769 ^ w973;
	assign w1036 = w1801 ^ w1004;
	assign w1002 = w1767 ^ w971;
	assign w1034 = w1799 ^ w1002;
	assign w1001 = w1766 ^ w970;
	assign w1033 = w1798 ^ w1001;
	assign w1069 = w1834 ^ w1037;
	assign w22853 = w1069 ^ w1063;
	assign w1068 = w1833 ^ w1036;
	assign w1066 = w1831 ^ w1034;
	assign w22766 = w1066 ^ w1068;
	assign w22852 = w1066 ^ w1069;
	assign w1065 = w1830 ^ w1033;
	assign w22763 = w1063 ^ w1065;
	assign w22844 = w22763 ^ w22852;
	assign w44332 = w22937 ^ w22939;
	assign w22895 = w44332 ^ w22892;
	assign w22992 = w22894 ^ w22895;
	assign w48093 = ~w22992;
	assign w967 = w1732 ^ w48093;
	assign w998 = w1763 ^ w967;
	assign w1030 = w1795 ^ w998;
	assign w1062 = w1827 ^ w1030;
	assign w22770 = w1062 ^ w1068;
	assign w22843 = w1062 ^ w22844;
	assign w22882 = w22886 ^ w44332;
	assign w22885 = w22924 ^ w22882;
	assign w22989 = w22884 ^ w22885;
	assign w22881 = w22905 ^ w22882;
	assign w48095 = w22880 ^ w22881;
	assign w48098 = ~w22989;
	assign w972 = w1737 ^ w48098;
	assign w969 = w1734 ^ w48095;
	assign w1003 = w1768 ^ w972;
	assign w1035 = w1800 ^ w1003;
	assign w1000 = w1765 ^ w969;
	assign w1032 = w1797 ^ w1000;
	assign w1067 = w1832 ^ w1035;
	assign w22764 = w1067 ^ w1069;
	assign w22847 = w22764 ^ w22770;
	assign w22850 = w1067 ^ w22770;
	assign w22846 = w1063 ^ w22850;
	assign w22726 = w22766 ^ w22764;
	assign w22842 = w22763 ^ w22726;
	assign w22725 = w22766 ^ w1067;
	assign w22849 = w1062 ^ w22725;
	assign w22835 = w22849 & w1062;
	assign w22833 = w22850 & w22846;
	assign w1064 = w1829 ^ w1032;
	assign w22765 = w1064 ^ w22763;
	assign w22841 = w1068 ^ w22765;
	assign w22838 = w1067 ^ w22765;
	assign w22840 = w22770 ^ w22765;
	assign w22780 = w1063 ^ w1064;
	assign w22845 = w22780 ^ w22847;
	assign w22848 = w22852 ^ w22780;
	assign w22854 = w1064 ^ w1066;
	assign w22839 = w22764 ^ w22854;
	assign w22740 = w1065 ^ w1064;
	assign w22851 = w1069 ^ w1064;
	assign w22837 = w22844 & w22848;
	assign w22769 = w22837 ^ w22766;
	assign w22836 = w22845 & w22843;
	assign w22834 = w22853 & w22838;
	assign w22768 = w22834 ^ w22764;
	assign w22832 = w22847 & w22840;
	assign w22831 = w22852 & w22841;
	assign w22767 = w22831 ^ w22765;
	assign w22773 = w22769 ^ w22767;
	assign w22778 = w1069 ^ w22773;
	assign w22830 = w22854 & w22839;
	assign w22787 = w22830 ^ w22836;
	assign w22828 = w22787 ^ w22778;
	assign w22739 = w22830 ^ w22831;
	assign w22786 = w22739 ^ w22740;
	assign w22785 = w22786 ^ w22768;
	assign w22827 = w22833 ^ w22785;
	assign w22829 = w22851 & w22842;
	assign w22824 = w22828 & w22827;
	assign w44323 = w22829 ^ w22832;
	assign w22742 = w22768 ^ w44323;
	assign w22826 = w22742 ^ w22767;
	assign w22823 = w22824 ^ w22826;
	assign w22782 = w22830 ^ w44323;
	assign w22738 = w22833 ^ w22782;
	assign w22820 = w1063 ^ w22738;
	assign w44326 = w22829 ^ w22835;
	assign w22741 = w22773 ^ w44326;
	assign w22784 = w1067 ^ w22741;
	assign w22819 = w22824 ^ w22784;
	assign w22818 = w22819 & w22820;
	assign w22816 = w22824 ^ w22818;
	assign w22737 = w22818 ^ w22782;
	assign w22736 = w22818 ^ w22835;
	assign w22731 = w22736 ^ w22832;
	assign w22815 = w22826 & w22816;
	assign w22813 = w22815 ^ w22823;
	assign w44325 = w22815 ^ w22833;
	assign w22807 = w44325 ^ w22785;
	assign w22796 = w22807 & w22848;
	assign w22805 = w22807 & w22844;
	assign w22774 = w1063 ^ w44325;
	assign w22814 = w22774 ^ w22737;
	assign w22804 = w22814 & w22843;
	assign w22795 = w22814 & w22845;
	assign w22817 = w22818 ^ w22826;
	assign w22803 = w22817 & w1062;
	assign w22794 = w22817 & w22849;
	assign w22779 = w44326 ^ w22764;
	assign w22825 = w22787 ^ w22779;
	assign w22822 = w22825 & w22823;
	assign w22821 = w22822 ^ w22784;
	assign w22733 = w22822 ^ w22834;
	assign w22729 = w22733 ^ w22769;
	assign w22732 = w1069 ^ w22729;
	assign w22809 = w22731 ^ w22732;
	assign w22730 = w22822 ^ w22778;
	assign w22728 = w1067 ^ w22729;
	assign w22812 = w22821 & w22813;
	assign w22777 = w22812 ^ w22787;
	assign w22811 = w22777 ^ w22779;
	assign w22735 = w22812 ^ w22836;
	assign w22727 = w22774 ^ w22735;
	assign w22734 = w22764 ^ w22727;
	assign w22810 = w22731 ^ w22734;
	assign w22808 = w22777 ^ w22730;
	assign w22806 = w22727 ^ w22728;
	assign w22802 = w22808 & w22838;
	assign w22801 = w22811 & w22850;
	assign w22800 = w22821 & w22840;
	assign w22744 = w22800 ^ w22801;
	assign w22799 = w22809 & w22841;
	assign w22798 = w22806 & w22839;
	assign w22759 = w22798 ^ w22801;
	assign w22756 = ~w22759;
	assign w22755 = w22798 ^ w22799;
	assign w22797 = w22810 & w22842;
	assign w22793 = w22808 & w22853;
	assign w22775 = w22793 ^ w22797;
	assign w22760 = w22802 ^ w22793;
	assign w22753 = ~w22775;
	assign w22792 = w22811 & w22846;
	assign w22762 = w22800 ^ w22792;
	assign w22791 = w22821 & w22847;
	assign w22752 = w22753 ^ w22791;
	assign w22790 = w22809 & w22852;
	assign w22789 = w22806 & w22854;
	assign w22788 = w22810 & w22851;
	assign w22754 = w22799 ^ w22788;
	assign w22750 = ~w22754;
	assign w44324 = w22789 ^ w22790;
	assign w22771 = w22795 ^ w44324;
	assign w22772 = w22796 ^ w22771;
	assign w22776 = w22804 ^ w22772;
	assign w22745 = w22803 ^ w22776;
	assign w48128 = w22744 ^ w22745;
	assign w1097 = w1862 ^ w48128;
	assign w1129 = w874 ^ w1097;
	assign w1161 = w906 ^ w1129;
	assign w1193 = w938 ^ w1161;
	assign w22781 = w22805 ^ w22776;
	assign w22856 = w22781 ^ w22755;
	assign w48131 = ~w22856;
	assign w1100 = w1865 ^ w48131;
	assign w1132 = w877 ^ w1100;
	assign w1164 = w909 ^ w1132;
	assign w1196 = w941 ^ w1164;
	assign w22758 = w22762 ^ w44324;
	assign w22757 = w22753 ^ w22758;
	assign w22857 = w22756 ^ w22757;
	assign w48126 = ~w22857;
	assign w1095 = w1860 ^ w48126;
	assign w1127 = w872 ^ w1095;
	assign w1159 = w904 ^ w1127;
	assign w1191 = w936 ^ w1159;
	assign w34957 = w1191 ^ w1193;
	assign w44327 = w22801 ^ w22802;
	assign w48129 = w44327 ^ w22781;
	assign w1098 = w1863 ^ w48129;
	assign w1130 = w875 ^ w1098;
	assign w1162 = w907 ^ w1130;
	assign w1194 = w939 ^ w1162;
	assign w34960 = w1194 ^ w1196;
	assign w22783 = w22798 ^ w44327;
	assign w22749 = w22794 ^ w22783;
	assign w22746 = ~w22749;
	assign w22743 = w22799 ^ w22783;
	assign w48132 = w22772 ^ w22743;
	assign w1101 = w1866 ^ w48132;
	assign w1133 = w878 ^ w1101;
	assign w1165 = w910 ^ w1133;
	assign w1197 = w942 ^ w1165;
	assign w35046 = w1194 ^ w1197;
	assign w35038 = w34957 ^ w35046;
	assign w35047 = w1197 ^ w1191;
	assign w44328 = w22803 ^ w22805;
	assign w22761 = w44328 ^ w22758;
	assign w22858 = w22760 ^ w22761;
	assign w48125 = ~w22858;
	assign w1094 = w1859 ^ w48125;
	assign w1126 = w871 ^ w1094;
	assign w1158 = w903 ^ w1126;
	assign w1190 = w935 ^ w1158;
	assign w34964 = w1190 ^ w1196;
	assign w35037 = w1190 ^ w35038;
	assign w22748 = w22752 ^ w44328;
	assign w22751 = w22790 ^ w22748;
	assign w22855 = w22750 ^ w22751;
	assign w22747 = w22771 ^ w22748;
	assign w48127 = w22746 ^ w22747;
	assign w48130 = ~w22855;
	assign w1099 = w1864 ^ w48130;
	assign w1131 = w876 ^ w1099;
	assign w1096 = w1861 ^ w48127;
	assign w1128 = w873 ^ w1096;
	assign w1163 = w908 ^ w1131;
	assign w1160 = w905 ^ w1128;
	assign w1192 = w937 ^ w1160;
	assign w34959 = w1192 ^ w34957;
	assign w35035 = w1196 ^ w34959;
	assign w35034 = w34964 ^ w34959;
	assign w34974 = w1191 ^ w1192;
	assign w35042 = w35046 ^ w34974;
	assign w35048 = w1192 ^ w1194;
	assign w34934 = w1193 ^ w1192;
	assign w35045 = w1197 ^ w1192;
	assign w35031 = w35038 & w35042;
	assign w34963 = w35031 ^ w34960;
	assign w35025 = w35046 & w35035;
	assign w34961 = w35025 ^ w34959;
	assign w34967 = w34963 ^ w34961;
	assign w34972 = w1197 ^ w34967;
	assign w1195 = w940 ^ w1163;
	assign w35032 = w1195 ^ w34959;
	assign w34958 = w1195 ^ w1197;
	assign w35033 = w34958 ^ w35048;
	assign w35041 = w34958 ^ w34964;
	assign w35039 = w34974 ^ w35041;
	assign w35044 = w1195 ^ w34964;
	assign w35040 = w1191 ^ w35044;
	assign w34920 = w34960 ^ w34958;
	assign w35036 = w34957 ^ w34920;
	assign w34919 = w34960 ^ w1195;
	assign w35043 = w1190 ^ w34919;
	assign w35030 = w35039 & w35037;
	assign w35029 = w35043 & w1190;
	assign w35028 = w35047 & w35032;
	assign w34962 = w35028 ^ w34958;
	assign w35027 = w35044 & w35040;
	assign w35026 = w35041 & w35034;
	assign w35024 = w35048 & w35033;
	assign w34981 = w35024 ^ w35030;
	assign w35022 = w34981 ^ w34972;
	assign w34933 = w35024 ^ w35025;
	assign w34980 = w34933 ^ w34934;
	assign w34979 = w34980 ^ w34962;
	assign w35021 = w35027 ^ w34979;
	assign w35023 = w35045 & w35036;
	assign w35018 = w35022 & w35021;
	assign w44834 = w35023 ^ w35029;
	assign w34935 = w34967 ^ w44834;
	assign w34978 = w1195 ^ w34935;
	assign w35013 = w35018 ^ w34978;
	assign w34973 = w44834 ^ w34958;
	assign w35019 = w34981 ^ w34973;
	assign w44835 = w35023 ^ w35026;
	assign w34976 = w35024 ^ w44835;
	assign w34932 = w35027 ^ w34976;
	assign w35014 = w1191 ^ w34932;
	assign w35012 = w35013 & w35014;
	assign w34931 = w35012 ^ w34976;
	assign w35010 = w35018 ^ w35012;
	assign w34930 = w35012 ^ w35029;
	assign w34925 = w34930 ^ w35026;
	assign w34936 = w34962 ^ w44835;
	assign w35020 = w34936 ^ w34961;
	assign w35011 = w35012 ^ w35020;
	assign w35017 = w35018 ^ w35020;
	assign w35016 = w35019 & w35017;
	assign w35015 = w35016 ^ w34978;
	assign w34927 = w35016 ^ w35028;
	assign w34923 = w34927 ^ w34963;
	assign w34926 = w1197 ^ w34923;
	assign w35003 = w34925 ^ w34926;
	assign w34924 = w35016 ^ w34972;
	assign w34922 = w1195 ^ w34923;
	assign w35009 = w35020 & w35010;
	assign w35007 = w35009 ^ w35017;
	assign w35006 = w35015 & w35007;
	assign w34971 = w35006 ^ w34981;
	assign w35005 = w34971 ^ w34973;
	assign w34929 = w35006 ^ w35030;
	assign w35002 = w34971 ^ w34924;
	assign w34997 = w35011 & w1190;
	assign w34996 = w35002 & w35032;
	assign w34995 = w35005 & w35044;
	assign w34994 = w35015 & w35034;
	assign w34938 = w34994 ^ w34995;
	assign w34993 = w35003 & w35035;
	assign w34988 = w35011 & w35043;
	assign w34987 = w35002 & w35047;
	assign w34954 = w34996 ^ w34987;
	assign w34986 = w35005 & w35040;
	assign w34956 = w34994 ^ w34986;
	assign w34985 = w35015 & w35041;
	assign w34984 = w35003 & w35046;
	assign w44837 = w34995 ^ w34996;
	assign w44839 = w35009 ^ w35027;
	assign w35001 = w44839 ^ w34979;
	assign w34999 = w35001 & w35038;
	assign w44838 = w34997 ^ w34999;
	assign w34990 = w35001 & w35042;
	assign w34968 = w1191 ^ w44839;
	assign w35008 = w34968 ^ w34931;
	assign w34921 = w34968 ^ w34929;
	assign w34928 = w34958 ^ w34921;
	assign w35004 = w34925 ^ w34928;
	assign w35000 = w34921 ^ w34922;
	assign w34998 = w35008 & w35037;
	assign w34992 = w35000 & w35033;
	assign w34977 = w34992 ^ w44837;
	assign w34953 = w34992 ^ w34995;
	assign w34950 = ~w34953;
	assign w34949 = w34992 ^ w34993;
	assign w34943 = w34988 ^ w34977;
	assign w34940 = ~w34943;
	assign w34937 = w34993 ^ w34977;
	assign w34991 = w35004 & w35036;
	assign w34969 = w34987 ^ w34991;
	assign w34947 = ~w34969;
	assign w34946 = w34947 ^ w34985;
	assign w34942 = w34946 ^ w44838;
	assign w34945 = w34984 ^ w34942;
	assign w34989 = w35008 & w35039;
	assign w34983 = w35000 & w35048;
	assign w34982 = w35004 & w35045;
	assign w34948 = w34993 ^ w34982;
	assign w34944 = ~w34948;
	assign w35049 = w34944 ^ w34945;
	assign w48170 = ~w35049;
	assign w1235 = w980 ^ w48170;
	assign w1266 = w1011 ^ w1235;
	assign w1298 = w1043 ^ w1266;
	assign w1330 = w1075 ^ w1298;
	assign w44836 = w34983 ^ w34984;
	assign w34965 = w34989 ^ w44836;
	assign w34966 = w34990 ^ w34965;
	assign w48172 = w34966 ^ w34937;
	assign w34970 = w34998 ^ w34966;
	assign w34975 = w34999 ^ w34970;
	assign w48169 = w44837 ^ w34975;
	assign w35050 = w34975 ^ w34949;
	assign w48171 = ~w35050;
	assign w34941 = w34965 ^ w34942;
	assign w1234 = w979 ^ w48169;
	assign w1265 = w1010 ^ w1234;
	assign w1297 = w1042 ^ w1265;
	assign w1329 = w1074 ^ w1297;
	assign w1237 = w982 ^ w48172;
	assign w1268 = w1013 ^ w1237;
	assign w48167 = w34940 ^ w34941;
	assign w1232 = w977 ^ w48167;
	assign w1263 = w1008 ^ w1232;
	assign w1295 = w1040 ^ w1263;
	assign w34939 = w34997 ^ w34970;
	assign w1327 = w1072 ^ w1295;
	assign w34914 = w1327 ^ w1329;
	assign w1236 = w981 ^ w48171;
	assign w1267 = w1012 ^ w1236;
	assign w1299 = w1044 ^ w1267;
	assign w1331 = w1076 ^ w1299;
	assign w34826 = w1329 ^ w1331;
	assign w34785 = w34826 ^ w1330;
	assign w48168 = w34938 ^ w34939;
	assign w1233 = w978 ^ w48168;
	assign w1264 = w1009 ^ w1233;
	assign w1296 = w1041 ^ w1264;
	assign w1328 = w1073 ^ w1296;
	assign w34800 = w1328 ^ w1327;
	assign w34952 = w34956 ^ w44836;
	assign w34955 = w44838 ^ w34952;
	assign w35052 = w34954 ^ w34955;
	assign w34951 = w34947 ^ w34952;
	assign w35051 = w34950 ^ w34951;
	assign w48165 = ~w35052;
	assign w48166 = ~w35051;
	assign w1231 = w976 ^ w48166;
	assign w1262 = w1007 ^ w1231;
	assign w1294 = w1039 ^ w1262;
	assign w1230 = w975 ^ w48165;
	assign w1261 = w1006 ^ w1230;
	assign w1293 = w1038 ^ w1261;
	assign w1326 = w1071 ^ w1294;
	assign w34823 = w1326 ^ w1328;
	assign w34825 = w1327 ^ w34823;
	assign w34901 = w1331 ^ w34825;
	assign w34898 = w1330 ^ w34825;
	assign w34840 = w1326 ^ w1327;
	assign w1325 = w1070 ^ w1293;
	assign w34830 = w1325 ^ w1331;
	assign w34900 = w34830 ^ w34825;
	assign w34910 = w1330 ^ w34830;
	assign w34906 = w1326 ^ w34910;
	assign w34909 = w1325 ^ w34785;
	assign w34895 = w34909 & w1325;
	assign w34893 = w34910 & w34906;
	assign w1300 = w1045 ^ w1268;
	assign w1332 = w1077 ^ w1300;
	assign w34824 = w1330 ^ w1332;
	assign w34899 = w34824 ^ w34914;
	assign w34912 = w1329 ^ w1332;
	assign w34908 = w34912 ^ w34840;
	assign w34907 = w34824 ^ w34830;
	assign w34905 = w34840 ^ w34907;
	assign w34904 = w34823 ^ w34912;
	assign w34903 = w1325 ^ w34904;
	assign w34786 = w34826 ^ w34824;
	assign w34902 = w34823 ^ w34786;
	assign w34913 = w1332 ^ w1326;
	assign w34911 = w1332 ^ w1327;
	assign w34897 = w34904 & w34908;
	assign w34829 = w34897 ^ w34826;
	assign w34896 = w34905 & w34903;
	assign w34894 = w34913 & w34898;
	assign w34828 = w34894 ^ w34824;
	assign w34892 = w34907 & w34900;
	assign w34891 = w34912 & w34901;
	assign w34827 = w34891 ^ w34825;
	assign w34833 = w34829 ^ w34827;
	assign w34838 = w1332 ^ w34833;
	assign w34890 = w34914 & w34899;
	assign w34847 = w34890 ^ w34896;
	assign w34888 = w34847 ^ w34838;
	assign w34799 = w34890 ^ w34891;
	assign w34846 = w34799 ^ w34800;
	assign w34845 = w34846 ^ w34828;
	assign w34887 = w34893 ^ w34845;
	assign w34889 = w34911 & w34902;
	assign w34884 = w34888 & w34887;
	assign w44829 = w34889 ^ w34895;
	assign w34839 = w44829 ^ w34824;
	assign w34885 = w34847 ^ w34839;
	assign w34801 = w34833 ^ w44829;
	assign w34844 = w1330 ^ w34801;
	assign w34879 = w34884 ^ w34844;
	assign w44830 = w34889 ^ w34892;
	assign w34842 = w34890 ^ w44830;
	assign w34798 = w34893 ^ w34842;
	assign w34880 = w1326 ^ w34798;
	assign w34878 = w34879 & w34880;
	assign w34797 = w34878 ^ w34842;
	assign w34796 = w34878 ^ w34895;
	assign w34791 = w34796 ^ w34892;
	assign w34876 = w34884 ^ w34878;
	assign w34802 = w34828 ^ w44830;
	assign w34886 = w34802 ^ w34827;
	assign w34877 = w34878 ^ w34886;
	assign w34883 = w34884 ^ w34886;
	assign w34882 = w34885 & w34883;
	assign w34881 = w34882 ^ w34844;
	assign w34793 = w34882 ^ w34894;
	assign w34789 = w34793 ^ w34829;
	assign w34792 = w1332 ^ w34789;
	assign w34869 = w34791 ^ w34792;
	assign w34790 = w34882 ^ w34838;
	assign w34788 = w1330 ^ w34789;
	assign w34875 = w34886 & w34876;
	assign w34873 = w34875 ^ w34883;
	assign w34872 = w34881 & w34873;
	assign w34837 = w34872 ^ w34847;
	assign w34871 = w34837 ^ w34839;
	assign w34795 = w34872 ^ w34896;
	assign w34868 = w34837 ^ w34790;
	assign w34863 = w34877 & w1325;
	assign w34862 = w34868 & w34898;
	assign w34861 = w34871 & w34910;
	assign w34860 = w34881 & w34900;
	assign w34804 = w34860 ^ w34861;
	assign w34859 = w34869 & w34901;
	assign w34854 = w34877 & w34909;
	assign w34853 = w34868 & w34913;
	assign w34820 = w34862 ^ w34853;
	assign w34852 = w34871 & w34906;
	assign w34822 = w34860 ^ w34852;
	assign w34851 = w34881 & w34907;
	assign w34850 = w34869 & w34912;
	assign w44831 = w34861 ^ w34862;
	assign w44833 = w34875 ^ w34893;
	assign w34834 = w1326 ^ w44833;
	assign w34874 = w34834 ^ w34797;
	assign w34855 = w34874 & w34905;
	assign w34864 = w34874 & w34903;
	assign w34787 = w34834 ^ w34795;
	assign w34794 = w34824 ^ w34787;
	assign w34870 = w34791 ^ w34794;
	assign w34857 = w34870 & w34902;
	assign w34835 = w34853 ^ w34857;
	assign w34813 = ~w34835;
	assign w34812 = w34813 ^ w34851;
	assign w34866 = w34787 ^ w34788;
	assign w34849 = w34866 & w34914;
	assign w34848 = w34870 & w34911;
	assign w34814 = w34859 ^ w34848;
	assign w34810 = ~w34814;
	assign w43596 = w34849 ^ w34850;
	assign w34818 = w34822 ^ w43596;
	assign w34817 = w34813 ^ w34818;
	assign w34831 = w34855 ^ w43596;
	assign w34858 = w34866 & w34899;
	assign w34815 = w34858 ^ w34859;
	assign w34843 = w34858 ^ w44831;
	assign w34809 = w34854 ^ w34843;
	assign w34806 = ~w34809;
	assign w34803 = w34859 ^ w34843;
	assign w34819 = w34858 ^ w34861;
	assign w34816 = ~w34819;
	assign w34917 = w34816 ^ w34817;
	assign w48198 = ~w34917;
	assign w1358 = w1103 ^ w48198;
	assign w401 = w1135 ^ w1358;
	assign w433 = w1167 ^ w401;
	assign w465 = w1199 ^ w433;
	assign w34867 = w44833 ^ w34845;
	assign w34865 = w34867 & w34904;
	assign w34856 = w34867 & w34908;
	assign w34832 = w34856 ^ w34831;
	assign w34836 = w34864 ^ w34832;
	assign w34841 = w34865 ^ w34836;
	assign w48201 = w44831 ^ w34841;
	assign w34916 = w34841 ^ w34815;
	assign w34805 = w34863 ^ w34836;
	assign w48200 = w34804 ^ w34805;
	assign w48204 = w34832 ^ w34803;
	assign w48203 = ~w34916;
	assign w1360 = w1105 ^ w48200;
	assign w403 = w1137 ^ w1360;
	assign w1363 = w1108 ^ w48203;
	assign w406 = w1140 ^ w1363;
	assign w1364 = w1109 ^ w48204;
	assign w1361 = w1106 ^ w48201;
	assign w404 = w1138 ^ w1361;
	assign w436 = w1170 ^ w404;
	assign w468 = w1202 ^ w436;
	assign w435 = w1169 ^ w403;
	assign w467 = w1201 ^ w435;
	assign w37503 = w465 ^ w467;
	assign w44832 = w34863 ^ w34865;
	assign w34821 = w44832 ^ w34818;
	assign w34918 = w34820 ^ w34821;
	assign w48197 = ~w34918;
	assign w1357 = w1102 ^ w48197;
	assign w400 = w1134 ^ w1357;
	assign w432 = w1166 ^ w400;
	assign w464 = w1198 ^ w432;
	assign w34808 = w34812 ^ w44832;
	assign w34811 = w34850 ^ w34808;
	assign w34915 = w34810 ^ w34811;
	assign w34807 = w34831 ^ w34808;
	assign w48199 = w34806 ^ w34807;
	assign w48202 = ~w34915;
	assign w1362 = w1107 ^ w48202;
	assign w1359 = w1104 ^ w48199;
	assign w402 = w1136 ^ w1359;
	assign w434 = w1168 ^ w402;
	assign w466 = w1200 ^ w434;
	assign w37505 = w466 ^ w37503;
	assign w37520 = w465 ^ w466;
	assign w37594 = w466 ^ w468;
	assign w37480 = w467 ^ w466;
	assign w405 = w1139 ^ w1362;
	assign w437 = w1171 ^ w405;
	assign w469 = w1203 ^ w437;
	assign w37578 = w469 ^ w37505;
	assign w407 = w1141 ^ w1364;
	assign w439 = w1173 ^ w407;
	assign w471 = w1205 ^ w439;
	assign w37504 = w469 ^ w471;
	assign w37579 = w37504 ^ w37594;
	assign w37592 = w468 ^ w471;
	assign w37588 = w37592 ^ w37520;
	assign w37584 = w37503 ^ w37592;
	assign w37583 = w464 ^ w37584;
	assign w37593 = w471 ^ w465;
	assign w37591 = w471 ^ w466;
	assign w37577 = w37584 & w37588;
	assign w37574 = w37593 & w37578;
	assign w37508 = w37574 ^ w37504;
	assign w37570 = w37594 & w37579;
	assign w438 = w1172 ^ w406;
	assign w470 = w1204 ^ w438;
	assign w37581 = w470 ^ w37505;
	assign w37506 = w468 ^ w470;
	assign w37509 = w37577 ^ w37506;
	assign w37510 = w464 ^ w470;
	assign w37580 = w37510 ^ w37505;
	assign w37587 = w37504 ^ w37510;
	assign w37585 = w37520 ^ w37587;
	assign w37590 = w469 ^ w37510;
	assign w37586 = w465 ^ w37590;
	assign w37466 = w37506 ^ w37504;
	assign w37582 = w37503 ^ w37466;
	assign w37465 = w37506 ^ w469;
	assign w37589 = w464 ^ w37465;
	assign w37576 = w37585 & w37583;
	assign w37527 = w37570 ^ w37576;
	assign w37575 = w37589 & w464;
	assign w37573 = w37590 & w37586;
	assign w37572 = w37587 & w37580;
	assign w37571 = w37592 & w37581;
	assign w37507 = w37571 ^ w37505;
	assign w37513 = w37509 ^ w37507;
	assign w37518 = w471 ^ w37513;
	assign w37568 = w37527 ^ w37518;
	assign w37479 = w37570 ^ w37571;
	assign w37526 = w37479 ^ w37480;
	assign w37525 = w37526 ^ w37508;
	assign w37567 = w37573 ^ w37525;
	assign w37569 = w37591 & w37582;
	assign w37564 = w37568 & w37567;
	assign w44942 = w37569 ^ w37572;
	assign w37482 = w37508 ^ w44942;
	assign w37566 = w37482 ^ w37507;
	assign w37563 = w37564 ^ w37566;
	assign w37522 = w37570 ^ w44942;
	assign w37478 = w37573 ^ w37522;
	assign w37560 = w465 ^ w37478;
	assign w44945 = w37569 ^ w37575;
	assign w37481 = w37513 ^ w44945;
	assign w37524 = w469 ^ w37481;
	assign w37559 = w37564 ^ w37524;
	assign w37558 = w37559 & w37560;
	assign w37556 = w37564 ^ w37558;
	assign w37477 = w37558 ^ w37522;
	assign w37476 = w37558 ^ w37575;
	assign w37471 = w37476 ^ w37572;
	assign w37555 = w37566 & w37556;
	assign w37553 = w37555 ^ w37563;
	assign w44944 = w37555 ^ w37573;
	assign w37547 = w44944 ^ w37525;
	assign w37536 = w37547 & w37588;
	assign w37545 = w37547 & w37584;
	assign w37514 = w465 ^ w44944;
	assign w37554 = w37514 ^ w37477;
	assign w37544 = w37554 & w37583;
	assign w37535 = w37554 & w37585;
	assign w37557 = w37558 ^ w37566;
	assign w37543 = w37557 & w464;
	assign w37534 = w37557 & w37589;
	assign w37519 = w44945 ^ w37504;
	assign w37565 = w37527 ^ w37519;
	assign w37562 = w37565 & w37563;
	assign w37561 = w37562 ^ w37524;
	assign w37473 = w37562 ^ w37574;
	assign w37469 = w37473 ^ w37509;
	assign w37472 = w471 ^ w37469;
	assign w37549 = w37471 ^ w37472;
	assign w37470 = w37562 ^ w37518;
	assign w37468 = w469 ^ w37469;
	assign w37552 = w37561 & w37553;
	assign w37517 = w37552 ^ w37527;
	assign w37551 = w37517 ^ w37519;
	assign w37475 = w37552 ^ w37576;
	assign w37467 = w37514 ^ w37475;
	assign w37474 = w37504 ^ w37467;
	assign w37550 = w37471 ^ w37474;
	assign w37548 = w37517 ^ w37470;
	assign w37546 = w37467 ^ w37468;
	assign w37542 = w37548 & w37578;
	assign w37541 = w37551 & w37590;
	assign w37540 = w37561 & w37580;
	assign w37484 = w37540 ^ w37541;
	assign w37539 = w37549 & w37581;
	assign w37538 = w37546 & w37579;
	assign w37499 = w37538 ^ w37541;
	assign w37496 = ~w37499;
	assign w37495 = w37538 ^ w37539;
	assign w37537 = w37550 & w37582;
	assign w37533 = w37548 & w37593;
	assign w37515 = w37533 ^ w37537;
	assign w37500 = w37542 ^ w37533;
	assign w37493 = ~w37515;
	assign w37532 = w37551 & w37586;
	assign w37502 = w37540 ^ w37532;
	assign w37531 = w37561 & w37587;
	assign w37492 = w37493 ^ w37531;
	assign w37530 = w37549 & w37592;
	assign w37529 = w37546 & w37594;
	assign w37528 = w37550 & w37591;
	assign w37494 = w37539 ^ w37528;
	assign w37490 = ~w37494;
	assign w44943 = w37529 ^ w37530;
	assign w37511 = w37535 ^ w44943;
	assign w37512 = w37536 ^ w37511;
	assign w37516 = w37544 ^ w37512;
	assign w37485 = w37543 ^ w37516;
	assign w48240 = w37484 ^ w37485;
	assign w37521 = w37545 ^ w37516;
	assign w37596 = w37521 ^ w37495;
	assign w48243 = ~w37596;
	assign w509 = w1243 ^ w48243;
	assign w541 = w1275 ^ w509;
	assign w573 = w1307 ^ w541;
	assign w605 = w1339 ^ w573;
	assign w37498 = w37502 ^ w44943;
	assign w37497 = w37493 ^ w37498;
	assign w37597 = w37496 ^ w37497;
	assign w48238 = ~w37597;
	assign w505 = w1239 ^ w48238;
	assign w536 = w1270 ^ w505;
	assign w568 = w1302 ^ w536;
	assign w600 = w1334 ^ w568;
	assign w44946 = w37541 ^ w37542;
	assign w48241 = w44946 ^ w37521;
	assign w37523 = w37538 ^ w44946;
	assign w37489 = w37534 ^ w37523;
	assign w37486 = ~w37489;
	assign w37483 = w37539 ^ w37523;
	assign w48244 = w37512 ^ w37483;
	assign w510 = w1244 ^ w48244;
	assign w542 = w1276 ^ w510;
	assign w574 = w1308 ^ w542;
	assign w606 = w1340 ^ w574;
	assign w38933 = w606 ^ w600;
	assign w44947 = w37543 ^ w37545;
	assign w37501 = w44947 ^ w37498;
	assign w37598 = w37500 ^ w37501;
	assign w48237 = ~w37598;
	assign w504 = w1238 ^ w48237;
	assign w535 = w1269 ^ w504;
	assign w567 = w1301 ^ w535;
	assign w599 = w1333 ^ w567;
	assign w38850 = w599 ^ w605;
	assign w37488 = w37492 ^ w44947;
	assign w37491 = w37530 ^ w37488;
	assign w37595 = w37490 ^ w37491;
	assign w37487 = w37511 ^ w37488;
	assign w48239 = w37486 ^ w37487;
	assign w48242 = ~w37595;
	assign w2047 = w1242 ^ w48242;
	assign w45168 = ~w2047;
	assign w540 = w1274 ^ w45168;
	assign w572 = w1306 ^ w540;
	assign w604 = w1338 ^ w572;
	assign w38844 = w604 ^ w606;
	assign w38927 = w38844 ^ w38850;
	assign w38930 = w604 ^ w38850;
	assign w38926 = w600 ^ w38930;
	assign w38913 = w38930 & w38926;
	assign w45169 = ~w2046;
	assign w1273 = w1018 ^ w45169;
	assign w1305 = w1050 ^ w1273;
	assign w1337 = w1082 ^ w1305;
	assign w37640 = w1337 ^ w1339;
	assign w37726 = w1337 ^ w1340;
	assign w37600 = w37640 ^ w37638;
	assign w37599 = w37640 ^ w1338;
	assign w37723 = w1333 ^ w37599;
	assign w37709 = w37723 & w1333;
	assign w508 = w45169 ^ w48241;
	assign w539 = w1273 ^ w508;
	assign w571 = w1305 ^ w539;
	assign w603 = w1337 ^ w571;
	assign w38846 = w603 ^ w605;
	assign w38932 = w603 ^ w606;
	assign w38806 = w38846 ^ w38844;
	assign w38805 = w38846 ^ w604;
	assign w38929 = w599 ^ w38805;
	assign w38915 = w599 & w38929;
	assign w45170 = ~w2045;
	assign w1017 = w1782 ^ w45170;
	assign w1049 = w1814 ^ w1017;
	assign w1081 = w1846 ^ w1049;
	assign w1241 = w45170 ^ w48176;
	assign w1272 = w1017 ^ w1241;
	assign w1304 = w1049 ^ w1272;
	assign w1336 = w1081 ^ w1304;
	assign w37637 = w1334 ^ w1336;
	assign w37718 = w37637 ^ w37726;
	assign w37717 = w1333 ^ w37718;
	assign w37716 = w37637 ^ w37600;
	assign w37905 = w1079 ^ w1081;
	assign w37986 = w37905 ^ w37994;
	assign w37985 = w1078 ^ w37986;
	assign w37984 = w37905 ^ w37868;
	assign w507 = w1241 ^ w48240;
	assign w538 = w1272 ^ w507;
	assign w570 = w1304 ^ w538;
	assign w602 = w1336 ^ w570;
	assign w38843 = w600 ^ w602;
	assign w38924 = w38843 ^ w38932;
	assign w38923 = w599 ^ w38924;
	assign w38922 = w38843 ^ w38806;
	assign w45171 = ~w2044;
	assign w1781 = w1526 ^ w45171;
	assign w1813 = w1558 ^ w1781;
	assign w1845 = w1590 ^ w1813;
	assign w985 = w45171 ^ w48111;
	assign w1016 = w1781 ^ w985;
	assign w1048 = w1813 ^ w1016;
	assign w1080 = w1845 ^ w1048;
	assign w37907 = w1080 ^ w37905;
	assign w37983 = w1084 ^ w37907;
	assign w37980 = w1083 ^ w37907;
	assign w37982 = w37912 ^ w37907;
	assign w37922 = w1079 ^ w1080;
	assign w37987 = w37922 ^ w37989;
	assign w37990 = w37994 ^ w37922;
	assign w37996 = w1080 ^ w1082;
	assign w37981 = w37906 ^ w37996;
	assign w37882 = w1081 ^ w1080;
	assign w37993 = w1085 ^ w1080;
	assign w37979 = w37986 & w37990;
	assign w37911 = w37979 ^ w37908;
	assign w37978 = w37987 & w37985;
	assign w37976 = w37995 & w37980;
	assign w37910 = w37976 ^ w37906;
	assign w37974 = w37989 & w37982;
	assign w37973 = w37994 & w37983;
	assign w37909 = w37973 ^ w37907;
	assign w37915 = w37911 ^ w37909;
	assign w37920 = w1085 ^ w37915;
	assign w37972 = w37996 & w37981;
	assign w37929 = w37972 ^ w37978;
	assign w37970 = w37929 ^ w37920;
	assign w37881 = w37972 ^ w37973;
	assign w37928 = w37881 ^ w37882;
	assign w37927 = w37928 ^ w37910;
	assign w37969 = w37975 ^ w37927;
	assign w37971 = w37993 & w37984;
	assign w37966 = w37970 & w37969;
	assign w38175 = w1845 ^ w38173;
	assign w38251 = w1849 ^ w38175;
	assign w38248 = w1848 ^ w38175;
	assign w38250 = w38180 ^ w38175;
	assign w38190 = w1844 ^ w1845;
	assign w38255 = w38190 ^ w38257;
	assign w38258 = w38262 ^ w38190;
	assign w38264 = w1845 ^ w1847;
	assign w38249 = w38174 ^ w38264;
	assign w38150 = w1846 ^ w1845;
	assign w38261 = w1850 ^ w1845;
	assign w38247 = w38254 & w38258;
	assign w38179 = w38247 ^ w38176;
	assign w38246 = w38255 & w38253;
	assign w38244 = w38263 & w38248;
	assign w38178 = w38244 ^ w38174;
	assign w38242 = w38257 & w38250;
	assign w38241 = w38262 & w38251;
	assign w38177 = w38241 ^ w38175;
	assign w38183 = w38179 ^ w38177;
	assign w38188 = w1850 ^ w38183;
	assign w38240 = w38264 & w38249;
	assign w38197 = w38240 ^ w38246;
	assign w38238 = w38197 ^ w38188;
	assign w38149 = w38240 ^ w38241;
	assign w38196 = w38149 ^ w38150;
	assign w38195 = w38196 ^ w38178;
	assign w38237 = w38243 ^ w38195;
	assign w38239 = w38261 & w38252;
	assign w38234 = w38238 & w38237;
	assign w1240 = w985 ^ w48175;
	assign w1271 = w1016 ^ w1240;
	assign w1303 = w1048 ^ w1271;
	assign w1335 = w1080 ^ w1303;
	assign w37639 = w1335 ^ w37637;
	assign w37715 = w1339 ^ w37639;
	assign w37712 = w1338 ^ w37639;
	assign w37714 = w37644 ^ w37639;
	assign w37654 = w1334 ^ w1335;
	assign w37719 = w37654 ^ w37721;
	assign w37722 = w37726 ^ w37654;
	assign w37728 = w1335 ^ w1337;
	assign w37713 = w37638 ^ w37728;
	assign w37614 = w1336 ^ w1335;
	assign w37725 = w1340 ^ w1335;
	assign w37711 = w37718 & w37722;
	assign w37643 = w37711 ^ w37640;
	assign w37710 = w37719 & w37717;
	assign w37708 = w37727 & w37712;
	assign w37642 = w37708 ^ w37638;
	assign w37706 = w37721 & w37714;
	assign w37705 = w37726 & w37715;
	assign w37641 = w37705 ^ w37639;
	assign w37647 = w37643 ^ w37641;
	assign w37652 = w1340 ^ w37647;
	assign w37704 = w37728 & w37713;
	assign w37661 = w37704 ^ w37710;
	assign w37702 = w37661 ^ w37652;
	assign w37613 = w37704 ^ w37705;
	assign w37660 = w37613 ^ w37614;
	assign w37659 = w37660 ^ w37642;
	assign w37701 = w37707 ^ w37659;
	assign w37703 = w37725 & w37716;
	assign w37698 = w37702 & w37701;
	assign w506 = w1240 ^ w48239;
	assign w537 = w1271 ^ w506;
	assign w569 = w1303 ^ w537;
	assign w601 = w1335 ^ w569;
	assign w38845 = w601 ^ w38843;
	assign w38921 = w605 ^ w38845;
	assign w38918 = w604 ^ w38845;
	assign w38920 = w38850 ^ w38845;
	assign w38860 = w600 ^ w601;
	assign w38925 = w38860 ^ w38927;
	assign w38928 = w38932 ^ w38860;
	assign w38934 = w601 ^ w603;
	assign w38919 = w38844 ^ w38934;
	assign w38820 = w602 ^ w601;
	assign w38931 = w606 ^ w601;
	assign w38917 = w38924 & w38928;
	assign w38849 = w38917 ^ w38846;
	assign w38916 = w38925 & w38923;
	assign w38914 = w38933 & w38918;
	assign w38848 = w38914 ^ w38844;
	assign w38912 = w38927 & w38920;
	assign w38911 = w38932 & w38921;
	assign w38847 = w38911 ^ w38845;
	assign w38853 = w38849 ^ w38847;
	assign w38858 = w606 ^ w38853;
	assign w38910 = w38934 & w38919;
	assign w38867 = w38910 ^ w38916;
	assign w38908 = w38867 ^ w38858;
	assign w38819 = w38910 ^ w38911;
	assign w38866 = w38819 ^ w38820;
	assign w38865 = w38866 ^ w38848;
	assign w38907 = w38913 ^ w38865;
	assign w38909 = w38931 & w38922;
	assign w38904 = w38908 & w38907;
	assign w44948 = w37703 ^ w37709;
	assign w37653 = w44948 ^ w37638;
	assign w37699 = w37661 ^ w37653;
	assign w37615 = w37647 ^ w44948;
	assign w37658 = w1338 ^ w37615;
	assign w37693 = w37698 ^ w37658;
	assign w44949 = w37703 ^ w37706;
	assign w37656 = w37704 ^ w44949;
	assign w37612 = w37707 ^ w37656;
	assign w37694 = w1334 ^ w37612;
	assign w37692 = w37693 & w37694;
	assign w37690 = w37698 ^ w37692;
	assign w37611 = w37692 ^ w37656;
	assign w37610 = w37692 ^ w37709;
	assign w37605 = w37610 ^ w37706;
	assign w37616 = w37642 ^ w44949;
	assign w37700 = w37616 ^ w37641;
	assign w37691 = w37692 ^ w37700;
	assign w37697 = w37698 ^ w37700;
	assign w37696 = w37699 & w37697;
	assign w37695 = w37696 ^ w37658;
	assign w37607 = w37696 ^ w37708;
	assign w37603 = w37607 ^ w37643;
	assign w37606 = w1340 ^ w37603;
	assign w37683 = w37605 ^ w37606;
	assign w37604 = w37696 ^ w37652;
	assign w37602 = w1338 ^ w37603;
	assign w37689 = w37700 & w37690;
	assign w37687 = w37689 ^ w37697;
	assign w37686 = w37695 & w37687;
	assign w37651 = w37686 ^ w37661;
	assign w37685 = w37651 ^ w37653;
	assign w37609 = w37686 ^ w37710;
	assign w37682 = w37651 ^ w37604;
	assign w37677 = w37691 & w1333;
	assign w37676 = w37682 & w37712;
	assign w37675 = w37685 & w37724;
	assign w37674 = w37695 & w37714;
	assign w37618 = w37674 ^ w37675;
	assign w37673 = w37683 & w37715;
	assign w37668 = w37691 & w37723;
	assign w37667 = w37682 & w37727;
	assign w37634 = w37676 ^ w37667;
	assign w37666 = w37685 & w37720;
	assign w37636 = w37674 ^ w37666;
	assign w37665 = w37695 & w37721;
	assign w37664 = w37683 & w37726;
	assign w44950 = w37675 ^ w37676;
	assign w44952 = w37689 ^ w37707;
	assign w37648 = w1334 ^ w44952;
	assign w37688 = w37648 ^ w37611;
	assign w37601 = w37648 ^ w37609;
	assign w37608 = w37638 ^ w37601;
	assign w37684 = w37605 ^ w37608;
	assign w37680 = w37601 ^ w37602;
	assign w37678 = w37688 & w37717;
	assign w37672 = w37680 & w37713;
	assign w37633 = w37672 ^ w37675;
	assign w37630 = ~w37633;
	assign w37629 = w37672 ^ w37673;
	assign w37671 = w37684 & w37716;
	assign w37669 = w37688 & w37719;
	assign w37649 = w37667 ^ w37671;
	assign w37627 = ~w37649;
	assign w37626 = w37627 ^ w37665;
	assign w37663 = w37680 & w37728;
	assign w37662 = w37684 & w37725;
	assign w37628 = w37673 ^ w37662;
	assign w37624 = ~w37628;
	assign w43603 = w37663 ^ w37664;
	assign w37632 = w37636 ^ w43603;
	assign w37631 = w37627 ^ w37632;
	assign w37731 = w37630 ^ w37631;
	assign w48206 = ~w37731;
	assign w37645 = w37669 ^ w43603;
	assign w37657 = w37672 ^ w44950;
	assign w37623 = w37668 ^ w37657;
	assign w37620 = ~w37623;
	assign w37617 = w37673 ^ w37657;
	assign w37681 = w44952 ^ w37659;
	assign w37679 = w37681 & w37718;
	assign w37670 = w37681 & w37722;
	assign w37646 = w37670 ^ w37645;
	assign w37650 = w37678 ^ w37646;
	assign w37655 = w37679 ^ w37650;
	assign w48209 = w44950 ^ w37655;
	assign w37730 = w37655 ^ w37629;
	assign w37619 = w37677 ^ w37650;
	assign w48208 = w37618 ^ w37619;
	assign w48212 = w37646 ^ w37617;
	assign w48211 = ~w37730;
	assign w44951 = w37677 ^ w37679;
	assign w37635 = w44951 ^ w37632;
	assign w37732 = w37634 ^ w37635;
	assign w48205 = ~w37732;
	assign w37622 = w37626 ^ w44951;
	assign w37625 = w37664 ^ w37622;
	assign w37729 = w37624 ^ w37625;
	assign w37621 = w37645 ^ w37622;
	assign w48207 = w37620 ^ w37621;
	assign w48210 = ~w37729;
	assign w44959 = w37971 ^ w37974;
	assign w37884 = w37910 ^ w44959;
	assign w37968 = w37884 ^ w37909;
	assign w37965 = w37966 ^ w37968;
	assign w37924 = w37972 ^ w44959;
	assign w37880 = w37975 ^ w37924;
	assign w37962 = w1079 ^ w37880;
	assign w44962 = w37971 ^ w37977;
	assign w37883 = w37915 ^ w44962;
	assign w37926 = w1083 ^ w37883;
	assign w37961 = w37966 ^ w37926;
	assign w37960 = w37961 & w37962;
	assign w37959 = w37960 ^ w37968;
	assign w37958 = w37966 ^ w37960;
	assign w37879 = w37960 ^ w37924;
	assign w37878 = w37960 ^ w37977;
	assign w37873 = w37878 ^ w37974;
	assign w37957 = w37968 & w37958;
	assign w37955 = w37957 ^ w37965;
	assign w37945 = w37959 & w1078;
	assign w37936 = w37959 & w37991;
	assign w44961 = w37957 ^ w37975;
	assign w37949 = w44961 ^ w37927;
	assign w37947 = w37949 & w37986;
	assign w37938 = w37949 & w37990;
	assign w37916 = w1079 ^ w44961;
	assign w37956 = w37916 ^ w37879;
	assign w37946 = w37956 & w37985;
	assign w37937 = w37956 & w37987;
	assign w37921 = w44962 ^ w37906;
	assign w37967 = w37929 ^ w37921;
	assign w37964 = w37967 & w37965;
	assign w37963 = w37964 ^ w37926;
	assign w37875 = w37964 ^ w37976;
	assign w37871 = w37875 ^ w37911;
	assign w37874 = w1085 ^ w37871;
	assign w37951 = w37873 ^ w37874;
	assign w37872 = w37964 ^ w37920;
	assign w37870 = w1083 ^ w37871;
	assign w37954 = w37963 & w37955;
	assign w37919 = w37954 ^ w37929;
	assign w37953 = w37919 ^ w37921;
	assign w37877 = w37954 ^ w37978;
	assign w37869 = w37916 ^ w37877;
	assign w37876 = w37906 ^ w37869;
	assign w37952 = w37873 ^ w37876;
	assign w37950 = w37919 ^ w37872;
	assign w37948 = w37869 ^ w37870;
	assign w37944 = w37950 & w37980;
	assign w37943 = w37953 & w37992;
	assign w37942 = w37963 & w37982;
	assign w37886 = w37942 ^ w37943;
	assign w37941 = w37951 & w37983;
	assign w37940 = w37948 & w37981;
	assign w37901 = w37940 ^ w37943;
	assign w37898 = ~w37901;
	assign w37897 = w37940 ^ w37941;
	assign w37939 = w37952 & w37984;
	assign w37935 = w37950 & w37995;
	assign w37917 = w37935 ^ w37939;
	assign w37902 = w37944 ^ w37935;
	assign w37895 = ~w37917;
	assign w37934 = w37953 & w37988;
	assign w37904 = w37942 ^ w37934;
	assign w37933 = w37963 & w37989;
	assign w37894 = w37895 ^ w37933;
	assign w37932 = w37951 & w37994;
	assign w37931 = w37948 & w37996;
	assign w37930 = w37952 & w37993;
	assign w37896 = w37941 ^ w37930;
	assign w37892 = ~w37896;
	assign w44960 = w37931 ^ w37932;
	assign w37913 = w37937 ^ w44960;
	assign w37914 = w37938 ^ w37913;
	assign w37918 = w37946 ^ w37914;
	assign w37923 = w37947 ^ w37918;
	assign w37998 = w37923 ^ w37897;
	assign w37887 = w37945 ^ w37918;
	assign w48144 = w37886 ^ w37887;
	assign w48147 = ~w37998;
	assign w37900 = w37904 ^ w44960;
	assign w37899 = w37895 ^ w37900;
	assign w37999 = w37898 ^ w37899;
	assign w48142 = ~w37999;
	assign w44963 = w37943 ^ w37944;
	assign w48145 = w44963 ^ w37923;
	assign w37925 = w37940 ^ w44963;
	assign w37891 = w37936 ^ w37925;
	assign w37888 = ~w37891;
	assign w37885 = w37941 ^ w37925;
	assign w48148 = w37914 ^ w37885;
	assign w44964 = w37945 ^ w37947;
	assign w37903 = w44964 ^ w37900;
	assign w38000 = w37902 ^ w37903;
	assign w48141 = ~w38000;
	assign w37890 = w37894 ^ w44964;
	assign w37893 = w37932 ^ w37890;
	assign w37997 = w37892 ^ w37893;
	assign w37889 = w37913 ^ w37890;
	assign w48143 = w37888 ^ w37889;
	assign w48146 = ~w37997;
	assign w44970 = w38239 ^ w38245;
	assign w38151 = w38183 ^ w44970;
	assign w38194 = w1848 ^ w38151;
	assign w38229 = w38234 ^ w38194;
	assign w38189 = w44970 ^ w38174;
	assign w38235 = w38197 ^ w38189;
	assign w44971 = w38239 ^ w38242;
	assign w38192 = w38240 ^ w44971;
	assign w38148 = w38243 ^ w38192;
	assign w38230 = w1844 ^ w38148;
	assign w38228 = w38229 & w38230;
	assign w38226 = w38234 ^ w38228;
	assign w38146 = w38228 ^ w38245;
	assign w38141 = w38146 ^ w38242;
	assign w38147 = w38228 ^ w38192;
	assign w38152 = w38178 ^ w44971;
	assign w38236 = w38152 ^ w38177;
	assign w38227 = w38228 ^ w38236;
	assign w38233 = w38234 ^ w38236;
	assign w38232 = w38235 & w38233;
	assign w38231 = w38232 ^ w38194;
	assign w38143 = w38232 ^ w38244;
	assign w38139 = w38143 ^ w38179;
	assign w38142 = w1850 ^ w38139;
	assign w38219 = w38141 ^ w38142;
	assign w38140 = w38232 ^ w38188;
	assign w38138 = w1848 ^ w38139;
	assign w38225 = w38236 & w38226;
	assign w38223 = w38225 ^ w38233;
	assign w38222 = w38231 & w38223;
	assign w38187 = w38222 ^ w38197;
	assign w38221 = w38187 ^ w38189;
	assign w38145 = w38222 ^ w38246;
	assign w38218 = w38187 ^ w38140;
	assign w38213 = w38227 & w1843;
	assign w38212 = w38218 & w38248;
	assign w38211 = w38221 & w38260;
	assign w38210 = w38231 & w38250;
	assign w38154 = w38210 ^ w38211;
	assign w38209 = w38219 & w38251;
	assign w38204 = w38227 & w38259;
	assign w38203 = w38218 & w38263;
	assign w38170 = w38212 ^ w38203;
	assign w38202 = w38221 & w38256;
	assign w38172 = w38210 ^ w38202;
	assign w38201 = w38231 & w38257;
	assign w38200 = w38219 & w38262;
	assign w44973 = w38211 ^ w38212;
	assign w44975 = w38225 ^ w38243;
	assign w38217 = w44975 ^ w38195;
	assign w38206 = w38217 & w38258;
	assign w38215 = w38217 & w38254;
	assign w44974 = w38213 ^ w38215;
	assign w38184 = w1844 ^ w44975;
	assign w38224 = w38184 ^ w38147;
	assign w38137 = w38184 ^ w38145;
	assign w38144 = w38174 ^ w38137;
	assign w38220 = w38141 ^ w38144;
	assign w38216 = w38137 ^ w38138;
	assign w38214 = w38224 & w38253;
	assign w38208 = w38216 & w38249;
	assign w38193 = w38208 ^ w44973;
	assign w38169 = w38208 ^ w38211;
	assign w38166 = ~w38169;
	assign w38165 = w38208 ^ w38209;
	assign w38159 = w38204 ^ w38193;
	assign w38156 = ~w38159;
	assign w38153 = w38209 ^ w38193;
	assign w38207 = w38220 & w38252;
	assign w38185 = w38203 ^ w38207;
	assign w38163 = ~w38185;
	assign w38162 = w38163 ^ w38201;
	assign w38158 = w38162 ^ w44974;
	assign w38161 = w38200 ^ w38158;
	assign w38205 = w38224 & w38255;
	assign w38199 = w38216 & w38264;
	assign w38198 = w38220 & w38261;
	assign w38164 = w38209 ^ w38198;
	assign w38160 = ~w38164;
	assign w38265 = w38160 ^ w38161;
	assign w48082 = ~w38265;
	assign w1880 = w1625 ^ w48082;
	assign w892 = w1657 ^ w1880;
	assign w924 = w1689 ^ w892;
	assign w956 = w1721 ^ w924;
	assign w1115 = w1880 ^ w48146;
	assign w1147 = w892 ^ w1115;
	assign w1179 = w924 ^ w1147;
	assign w1370 = w1115 ^ w48210;
	assign w413 = w1147 ^ w1370;
	assign w445 = w1179 ^ w413;
	assign w1211 = w956 ^ w1179;
	assign w477 = w1211 ^ w445;
	assign w44972 = w38199 ^ w38200;
	assign w38181 = w38205 ^ w44972;
	assign w38157 = w38181 ^ w38158;
	assign w48079 = w38156 ^ w38157;
	assign w1877 = w1622 ^ w48079;
	assign w889 = w1654 ^ w1877;
	assign w921 = w1686 ^ w889;
	assign w953 = w1718 ^ w921;
	assign w1112 = w1877 ^ w48143;
	assign w1144 = w889 ^ w1112;
	assign w1176 = w921 ^ w1144;
	assign w1367 = w1112 ^ w48207;
	assign w410 = w1144 ^ w1367;
	assign w442 = w1176 ^ w410;
	assign w38182 = w38206 ^ w38181;
	assign w48084 = w38182 ^ w38153;
	assign w1882 = w1627 ^ w48084;
	assign w894 = w1659 ^ w1882;
	assign w926 = w1691 ^ w894;
	assign w958 = w1723 ^ w926;
	assign w1117 = w1882 ^ w48148;
	assign w1372 = w1117 ^ w48212;
	assign w1149 = w894 ^ w1117;
	assign w1181 = w926 ^ w1149;
	assign w36921 = w958 ^ w953;
	assign w36834 = w956 ^ w958;
	assign w38186 = w38214 ^ w38182;
	assign w38155 = w38213 ^ w38186;
	assign w48080 = w38154 ^ w38155;
	assign w1878 = w1623 ^ w48080;
	assign w1113 = w1878 ^ w48144;
	assign w890 = w1655 ^ w1878;
	assign w1145 = w890 ^ w1113;
	assign w922 = w1687 ^ w890;
	assign w1177 = w922 ^ w1145;
	assign w954 = w1719 ^ w922;
	assign w36810 = w954 ^ w953;
	assign w38191 = w38215 ^ w38186;
	assign w38266 = w38191 ^ w38165;
	assign w48083 = ~w38266;
	assign w1881 = w1626 ^ w48083;
	assign w893 = w1658 ^ w1881;
	assign w925 = w1690 ^ w893;
	assign w957 = w1722 ^ w925;
	assign w1116 = w1881 ^ w48147;
	assign w1148 = w893 ^ w1116;
	assign w1180 = w925 ^ w1148;
	assign w1371 = w1116 ^ w48211;
	assign w414 = w1148 ^ w1371;
	assign w446 = w1180 ^ w414;
	assign w48081 = w44973 ^ w38191;
	assign w1879 = w1624 ^ w48081;
	assign w1114 = w1879 ^ w48145;
	assign w1369 = w1114 ^ w48209;
	assign w1213 = w958 ^ w1181;
	assign w36566 = w1211 ^ w1213;
	assign w1212 = w957 ^ w1180;
	assign w478 = w1212 ^ w446;
	assign w1209 = w954 ^ w1177;
	assign w1208 = w953 ^ w1176;
	assign w36542 = w1209 ^ w1208;
	assign w36653 = w1213 ^ w1208;
	assign w474 = w1208 ^ w442;
	assign w415 = w1149 ^ w1372;
	assign w447 = w1181 ^ w415;
	assign w479 = w1213 ^ w447;
	assign w36298 = w477 ^ w479;
	assign w36385 = w479 ^ w474;
	assign w1368 = w1113 ^ w48208;
	assign w411 = w1145 ^ w1368;
	assign w443 = w1177 ^ w411;
	assign w475 = w1209 ^ w443;
	assign w36274 = w475 ^ w474;
	assign w891 = w1656 ^ w1879;
	assign w923 = w1688 ^ w891;
	assign w955 = w1720 ^ w923;
	assign w36836 = w955 ^ w957;
	assign w36922 = w955 ^ w958;
	assign w36924 = w953 ^ w955;
	assign w36909 = w36834 ^ w36924;
	assign w36796 = w36836 ^ w36834;
	assign w36795 = w36836 ^ w956;
	assign w36900 = w36924 & w36909;
	assign w1146 = w891 ^ w1114;
	assign w412 = w1146 ^ w1369;
	assign w1178 = w923 ^ w1146;
	assign w1210 = w955 ^ w1178;
	assign w36656 = w1208 ^ w1210;
	assign w36641 = w36566 ^ w36656;
	assign w36632 = w36656 & w36641;
	assign w444 = w1178 ^ w412;
	assign w476 = w1210 ^ w444;
	assign w36300 = w476 ^ w478;
	assign w36386 = w476 ^ w479;
	assign w36388 = w474 ^ w476;
	assign w36373 = w36298 ^ w36388;
	assign w36260 = w36300 ^ w36298;
	assign w36259 = w36300 ^ w477;
	assign w36364 = w36388 & w36373;
	assign w36568 = w1210 ^ w1212;
	assign w36527 = w36568 ^ w1211;
	assign w36654 = w1210 ^ w1213;
	assign w36528 = w36568 ^ w36566;
	assign w38168 = w38172 ^ w44972;
	assign w38171 = w44974 ^ w38168;
	assign w38268 = w38170 ^ w38171;
	assign w38167 = w38163 ^ w38168;
	assign w38267 = w38166 ^ w38167;
	assign w48077 = ~w38268;
	assign w1875 = w1620 ^ w48077;
	assign w887 = w1652 ^ w1875;
	assign w919 = w1684 ^ w887;
	assign w951 = w1716 ^ w919;
	assign w1110 = w1875 ^ w48141;
	assign w1142 = w887 ^ w1110;
	assign w36840 = w951 ^ w957;
	assign w36917 = w36834 ^ w36840;
	assign w36920 = w956 ^ w36840;
	assign w36919 = w951 ^ w36795;
	assign w36905 = w36919 & w951;
	assign w1365 = w1110 ^ w48205;
	assign w408 = w1142 ^ w1365;
	assign w48078 = ~w38267;
	assign w1876 = w1621 ^ w48078;
	assign w888 = w1653 ^ w1876;
	assign w920 = w1685 ^ w888;
	assign w952 = w1717 ^ w920;
	assign w1111 = w1876 ^ w48142;
	assign w1366 = w1111 ^ w48206;
	assign w1143 = w888 ^ w1111;
	assign w1175 = w920 ^ w1143;
	assign w409 = w1143 ^ w1366;
	assign w36833 = w952 ^ w954;
	assign w36835 = w953 ^ w36833;
	assign w36911 = w957 ^ w36835;
	assign w36908 = w956 ^ w36835;
	assign w36910 = w36840 ^ w36835;
	assign w36916 = w952 ^ w36920;
	assign w36914 = w36833 ^ w36922;
	assign w36913 = w951 ^ w36914;
	assign w36850 = w952 ^ w953;
	assign w36915 = w36850 ^ w36917;
	assign w36918 = w36922 ^ w36850;
	assign w36912 = w36833 ^ w36796;
	assign w36923 = w958 ^ w952;
	assign w36907 = w36914 & w36918;
	assign w36839 = w36907 ^ w36836;
	assign w36906 = w36915 & w36913;
	assign w36857 = w36900 ^ w36906;
	assign w36904 = w36923 & w36908;
	assign w36838 = w36904 ^ w36834;
	assign w36903 = w36920 & w36916;
	assign w36902 = w36917 & w36910;
	assign w36901 = w36922 & w36911;
	assign w36837 = w36901 ^ w36835;
	assign w36843 = w36839 ^ w36837;
	assign w36848 = w958 ^ w36843;
	assign w36898 = w36857 ^ w36848;
	assign w36809 = w36900 ^ w36901;
	assign w36856 = w36809 ^ w36810;
	assign w36855 = w36856 ^ w36838;
	assign w36897 = w36903 ^ w36855;
	assign w36899 = w36921 & w36912;
	assign w36894 = w36898 & w36897;
	assign w441 = w1175 ^ w409;
	assign w1174 = w919 ^ w1142;
	assign w440 = w1174 ^ w408;
	assign w1207 = w952 ^ w1175;
	assign w36565 = w1207 ^ w1209;
	assign w36567 = w1208 ^ w36565;
	assign w36643 = w1212 ^ w36567;
	assign w36640 = w1211 ^ w36567;
	assign w36646 = w36565 ^ w36654;
	assign w36582 = w1207 ^ w1208;
	assign w36650 = w36654 ^ w36582;
	assign w36644 = w36565 ^ w36528;
	assign w36655 = w1213 ^ w1207;
	assign w36639 = w36646 & w36650;
	assign w36571 = w36639 ^ w36568;
	assign w36636 = w36655 & w36640;
	assign w36570 = w36636 ^ w36566;
	assign w36633 = w36654 & w36643;
	assign w36569 = w36633 ^ w36567;
	assign w36575 = w36571 ^ w36569;
	assign w36580 = w1213 ^ w36575;
	assign w36541 = w36632 ^ w36633;
	assign w36588 = w36541 ^ w36542;
	assign w36587 = w36588 ^ w36570;
	assign w36631 = w36653 & w36644;
	assign w473 = w1207 ^ w441;
	assign w36297 = w473 ^ w475;
	assign w36299 = w474 ^ w36297;
	assign w36375 = w478 ^ w36299;
	assign w36372 = w477 ^ w36299;
	assign w36378 = w36297 ^ w36386;
	assign w36314 = w473 ^ w474;
	assign w36382 = w36386 ^ w36314;
	assign w36376 = w36297 ^ w36260;
	assign w36387 = w479 ^ w473;
	assign w36371 = w36378 & w36382;
	assign w36303 = w36371 ^ w36300;
	assign w36368 = w36387 & w36372;
	assign w36302 = w36368 ^ w36298;
	assign w36365 = w36386 & w36375;
	assign w36301 = w36365 ^ w36299;
	assign w36307 = w36303 ^ w36301;
	assign w36312 = w479 ^ w36307;
	assign w36273 = w36364 ^ w36365;
	assign w36320 = w36273 ^ w36274;
	assign w36319 = w36320 ^ w36302;
	assign w36363 = w36385 & w36376;
	assign w1206 = w951 ^ w1174;
	assign w36645 = w1206 ^ w36646;
	assign w36572 = w1206 ^ w1212;
	assign w36642 = w36572 ^ w36567;
	assign w36649 = w36566 ^ w36572;
	assign w36647 = w36582 ^ w36649;
	assign w36652 = w1211 ^ w36572;
	assign w36648 = w1207 ^ w36652;
	assign w36651 = w1206 ^ w36527;
	assign w36638 = w36647 & w36645;
	assign w36589 = w36632 ^ w36638;
	assign w36630 = w36589 ^ w36580;
	assign w36637 = w36651 & w1206;
	assign w36635 = w36652 & w36648;
	assign w36629 = w36635 ^ w36587;
	assign w36634 = w36649 & w36642;
	assign w36626 = w36630 & w36629;
	assign w472 = w1206 ^ w440;
	assign w36377 = w472 ^ w36378;
	assign w36304 = w472 ^ w478;
	assign w36374 = w36304 ^ w36299;
	assign w36381 = w36298 ^ w36304;
	assign w36379 = w36314 ^ w36381;
	assign w36384 = w477 ^ w36304;
	assign w36380 = w473 ^ w36384;
	assign w36383 = w472 ^ w36259;
	assign w36370 = w36379 & w36377;
	assign w36321 = w36364 ^ w36370;
	assign w36362 = w36321 ^ w36312;
	assign w36369 = w36383 & w472;
	assign w36367 = w36384 & w36380;
	assign w36361 = w36367 ^ w36319;
	assign w36366 = w36381 & w36374;
	assign w36358 = w36362 & w36361;
	assign w44891 = w36363 ^ w36366;
	assign w36276 = w36302 ^ w44891;
	assign w36360 = w36276 ^ w36301;
	assign w36357 = w36358 ^ w36360;
	assign w36316 = w36364 ^ w44891;
	assign w36272 = w36367 ^ w36316;
	assign w36354 = w473 ^ w36272;
	assign w44894 = w36363 ^ w36369;
	assign w36275 = w36307 ^ w44894;
	assign w36318 = w477 ^ w36275;
	assign w36353 = w36358 ^ w36318;
	assign w36352 = w36353 & w36354;
	assign w36351 = w36352 ^ w36360;
	assign w36350 = w36358 ^ w36352;
	assign w36271 = w36352 ^ w36316;
	assign w36270 = w36352 ^ w36369;
	assign w36265 = w36270 ^ w36366;
	assign w36349 = w36360 & w36350;
	assign w36347 = w36349 ^ w36357;
	assign w36337 = w36351 & w472;
	assign w36328 = w36351 & w36383;
	assign w44893 = w36349 ^ w36367;
	assign w36341 = w44893 ^ w36319;
	assign w36339 = w36341 & w36378;
	assign w36330 = w36341 & w36382;
	assign w36308 = w473 ^ w44893;
	assign w36348 = w36308 ^ w36271;
	assign w36338 = w36348 & w36377;
	assign w36329 = w36348 & w36379;
	assign w36313 = w44894 ^ w36298;
	assign w36359 = w36321 ^ w36313;
	assign w36356 = w36359 & w36357;
	assign w36355 = w36356 ^ w36318;
	assign w36267 = w36356 ^ w36368;
	assign w36263 = w36267 ^ w36303;
	assign w36266 = w479 ^ w36263;
	assign w36343 = w36265 ^ w36266;
	assign w36264 = w36356 ^ w36312;
	assign w36262 = w477 ^ w36263;
	assign w36346 = w36355 & w36347;
	assign w36311 = w36346 ^ w36321;
	assign w36345 = w36311 ^ w36313;
	assign w36269 = w36346 ^ w36370;
	assign w36261 = w36308 ^ w36269;
	assign w36268 = w36298 ^ w36261;
	assign w36344 = w36265 ^ w36268;
	assign w36342 = w36311 ^ w36264;
	assign w36340 = w36261 ^ w36262;
	assign w36336 = w36342 & w36372;
	assign w36335 = w36345 & w36384;
	assign w36334 = w36355 & w36374;
	assign w36278 = w36334 ^ w36335;
	assign w36333 = w36343 & w36375;
	assign w36332 = w36340 & w36373;
	assign w36293 = w36332 ^ w36335;
	assign w36290 = ~w36293;
	assign w36289 = w36332 ^ w36333;
	assign w36331 = w36344 & w36376;
	assign w36327 = w36342 & w36387;
	assign w36309 = w36327 ^ w36331;
	assign w36294 = w36336 ^ w36327;
	assign w36287 = ~w36309;
	assign w36326 = w36345 & w36380;
	assign w36296 = w36334 ^ w36326;
	assign w36325 = w36355 & w36381;
	assign w36286 = w36287 ^ w36325;
	assign w36324 = w36343 & w36386;
	assign w36323 = w36340 & w36388;
	assign w36322 = w36344 & w36385;
	assign w36288 = w36333 ^ w36322;
	assign w36284 = ~w36288;
	assign w44892 = w36323 ^ w36324;
	assign w36292 = w36296 ^ w44892;
	assign w36291 = w36287 ^ w36292;
	assign w36391 = w36290 ^ w36291;
	assign w48214 = ~w36391;
	assign w36305 = w36329 ^ w44892;
	assign w36306 = w36330 ^ w36305;
	assign w36310 = w36338 ^ w36306;
	assign w36315 = w36339 ^ w36310;
	assign w36390 = w36315 ^ w36289;
	assign w36279 = w36337 ^ w36310;
	assign w48216 = w36278 ^ w36279;
	assign w48219 = ~w36390;
	assign w44895 = w36335 ^ w36336;
	assign w48217 = w44895 ^ w36315;
	assign w36317 = w36332 ^ w44895;
	assign w36283 = w36328 ^ w36317;
	assign w36280 = ~w36283;
	assign w36277 = w36333 ^ w36317;
	assign w48220 = w36306 ^ w36277;
	assign w44896 = w36337 ^ w36339;
	assign w36295 = w44896 ^ w36292;
	assign w36392 = w36294 ^ w36295;
	assign w48213 = ~w36392;
	assign w36282 = w36286 ^ w44896;
	assign w36285 = w36324 ^ w36282;
	assign w36389 = w36284 ^ w36285;
	assign w36281 = w36305 ^ w36282;
	assign w48215 = w36280 ^ w36281;
	assign w48218 = ~w36389;
	assign w44902 = w36631 ^ w36637;
	assign w36543 = w36575 ^ w44902;
	assign w36586 = w1211 ^ w36543;
	assign w36621 = w36626 ^ w36586;
	assign w36581 = w44902 ^ w36566;
	assign w36627 = w36589 ^ w36581;
	assign w44903 = w36631 ^ w36634;
	assign w36584 = w36632 ^ w44903;
	assign w36540 = w36635 ^ w36584;
	assign w36622 = w1207 ^ w36540;
	assign w36620 = w36621 & w36622;
	assign w36538 = w36620 ^ w36637;
	assign w36618 = w36626 ^ w36620;
	assign w36539 = w36620 ^ w36584;
	assign w36533 = w36538 ^ w36634;
	assign w36544 = w36570 ^ w44903;
	assign w36628 = w36544 ^ w36569;
	assign w36619 = w36620 ^ w36628;
	assign w36625 = w36626 ^ w36628;
	assign w36624 = w36627 & w36625;
	assign w36623 = w36624 ^ w36586;
	assign w36535 = w36624 ^ w36636;
	assign w36531 = w36535 ^ w36571;
	assign w36534 = w1213 ^ w36531;
	assign w36611 = w36533 ^ w36534;
	assign w36532 = w36624 ^ w36580;
	assign w36530 = w1211 ^ w36531;
	assign w36617 = w36628 & w36618;
	assign w36615 = w36617 ^ w36625;
	assign w36614 = w36623 & w36615;
	assign w36579 = w36614 ^ w36589;
	assign w36613 = w36579 ^ w36581;
	assign w36537 = w36614 ^ w36638;
	assign w36610 = w36579 ^ w36532;
	assign w36605 = w36619 & w1206;
	assign w36604 = w36610 & w36640;
	assign w36603 = w36613 & w36652;
	assign w36602 = w36623 & w36642;
	assign w36546 = w36602 ^ w36603;
	assign w36601 = w36611 & w36643;
	assign w36596 = w36619 & w36651;
	assign w36595 = w36610 & w36655;
	assign w36562 = w36604 ^ w36595;
	assign w36594 = w36613 & w36648;
	assign w36564 = w36602 ^ w36594;
	assign w36593 = w36623 & w36649;
	assign w36592 = w36611 & w36654;
	assign w44905 = w36603 ^ w36604;
	assign w44907 = w36617 ^ w36635;
	assign w36609 = w44907 ^ w36587;
	assign w36607 = w36609 & w36646;
	assign w36598 = w36609 & w36650;
	assign w44906 = w36605 ^ w36607;
	assign w36576 = w1207 ^ w44907;
	assign w36616 = w36576 ^ w36539;
	assign w36529 = w36576 ^ w36537;
	assign w36536 = w36566 ^ w36529;
	assign w36612 = w36533 ^ w36536;
	assign w36608 = w36529 ^ w36530;
	assign w36606 = w36616 & w36645;
	assign w36600 = w36608 & w36641;
	assign w36585 = w36600 ^ w44905;
	assign w36561 = w36600 ^ w36603;
	assign w36558 = ~w36561;
	assign w36557 = w36600 ^ w36601;
	assign w36551 = w36596 ^ w36585;
	assign w36548 = ~w36551;
	assign w36545 = w36601 ^ w36585;
	assign w36599 = w36612 & w36644;
	assign w36577 = w36595 ^ w36599;
	assign w36555 = ~w36577;
	assign w36554 = w36555 ^ w36593;
	assign w36550 = w36554 ^ w44906;
	assign w36553 = w36592 ^ w36550;
	assign w36597 = w36616 & w36647;
	assign w36591 = w36608 & w36656;
	assign w36590 = w36612 & w36653;
	assign w36556 = w36601 ^ w36590;
	assign w36552 = ~w36556;
	assign w36657 = w36552 ^ w36553;
	assign w48154 = ~w36657;
	assign w44904 = w36591 ^ w36592;
	assign w36560 = w36564 ^ w44904;
	assign w36563 = w44906 ^ w36560;
	assign w36660 = w36562 ^ w36563;
	assign w36559 = w36555 ^ w36560;
	assign w36659 = w36558 ^ w36559;
	assign w48149 = ~w36660;
	assign w48150 = ~w36659;
	assign w36573 = w36597 ^ w44904;
	assign w36574 = w36598 ^ w36573;
	assign w36578 = w36606 ^ w36574;
	assign w36583 = w36607 ^ w36578;
	assign w48153 = w44905 ^ w36583;
	assign w36658 = w36583 ^ w36557;
	assign w36549 = w36573 ^ w36550;
	assign w48151 = w36548 ^ w36549;
	assign w36547 = w36605 ^ w36578;
	assign w48152 = w36546 ^ w36547;
	assign w48156 = w36574 ^ w36545;
	assign w48155 = ~w36658;
	assign w44914 = w36899 ^ w36905;
	assign w36849 = w44914 ^ w36834;
	assign w36895 = w36857 ^ w36849;
	assign w36811 = w36843 ^ w44914;
	assign w36854 = w956 ^ w36811;
	assign w36889 = w36894 ^ w36854;
	assign w44915 = w36899 ^ w36902;
	assign w36852 = w36900 ^ w44915;
	assign w36808 = w36903 ^ w36852;
	assign w36890 = w952 ^ w36808;
	assign w36888 = w36889 & w36890;
	assign w36886 = w36894 ^ w36888;
	assign w36807 = w36888 ^ w36852;
	assign w36806 = w36888 ^ w36905;
	assign w36801 = w36806 ^ w36902;
	assign w36812 = w36838 ^ w44915;
	assign w36896 = w36812 ^ w36837;
	assign w36887 = w36888 ^ w36896;
	assign w36893 = w36894 ^ w36896;
	assign w36892 = w36895 & w36893;
	assign w36891 = w36892 ^ w36854;
	assign w36803 = w36892 ^ w36904;
	assign w36799 = w36803 ^ w36839;
	assign w36802 = w958 ^ w36799;
	assign w36879 = w36801 ^ w36802;
	assign w36800 = w36892 ^ w36848;
	assign w36798 = w956 ^ w36799;
	assign w36885 = w36896 & w36886;
	assign w36883 = w36885 ^ w36893;
	assign w36882 = w36891 & w36883;
	assign w36847 = w36882 ^ w36857;
	assign w36881 = w36847 ^ w36849;
	assign w36805 = w36882 ^ w36906;
	assign w36878 = w36847 ^ w36800;
	assign w36873 = w36887 & w951;
	assign w36872 = w36878 & w36908;
	assign w36871 = w36881 & w36920;
	assign w36870 = w36891 & w36910;
	assign w36814 = w36870 ^ w36871;
	assign w36869 = w36879 & w36911;
	assign w36864 = w36887 & w36919;
	assign w36863 = w36878 & w36923;
	assign w36830 = w36872 ^ w36863;
	assign w36862 = w36881 & w36916;
	assign w36832 = w36870 ^ w36862;
	assign w36861 = w36891 & w36917;
	assign w36860 = w36879 & w36922;
	assign w44916 = w36871 ^ w36872;
	assign w44918 = w36885 ^ w36903;
	assign w36844 = w952 ^ w44918;
	assign w36884 = w36844 ^ w36807;
	assign w36874 = w36884 & w36913;
	assign w36865 = w36884 & w36915;
	assign w36797 = w36844 ^ w36805;
	assign w36876 = w36797 ^ w36798;
	assign w36868 = w36876 & w36909;
	assign w36829 = w36868 ^ w36871;
	assign w36826 = ~w36829;
	assign w36825 = w36868 ^ w36869;
	assign w36859 = w36876 & w36924;
	assign w43601 = w36859 ^ w36860;
	assign w36828 = w36832 ^ w43601;
	assign w36841 = w36865 ^ w43601;
	assign w36804 = w36834 ^ w36797;
	assign w36853 = w36868 ^ w44916;
	assign w36819 = w36864 ^ w36853;
	assign w36816 = ~w36819;
	assign w36813 = w36869 ^ w36853;
	assign w36880 = w36801 ^ w36804;
	assign w36858 = w36880 & w36921;
	assign w36824 = w36869 ^ w36858;
	assign w36820 = ~w36824;
	assign w36867 = w36880 & w36912;
	assign w36845 = w36863 ^ w36867;
	assign w36823 = ~w36845;
	assign w36827 = w36823 ^ w36828;
	assign w36927 = w36826 ^ w36827;
	assign w48086 = ~w36927;
	assign w960 = w1725 ^ w48086;
	assign w991 = w1756 ^ w960;
	assign w1023 = w1788 ^ w991;
	assign w1055 = w1820 ^ w1023;
	assign w36822 = w36823 ^ w36861;
	assign w1215 = w960 ^ w48150;
	assign w1246 = w991 ^ w1215;
	assign w1278 = w1023 ^ w1246;
	assign w1310 = w1055 ^ w1278;
	assign w481 = w1215 ^ w48214;
	assign w512 = w1246 ^ w481;
	assign w544 = w1278 ^ w512;
	assign w576 = w1310 ^ w544;
	assign w36877 = w44918 ^ w36855;
	assign w36875 = w36877 & w36914;
	assign w36866 = w36877 & w36918;
	assign w36842 = w36866 ^ w36841;
	assign w36846 = w36874 ^ w36842;
	assign w36851 = w36875 ^ w36846;
	assign w48089 = w44916 ^ w36851;
	assign w963 = w1728 ^ w48089;
	assign w994 = w1759 ^ w963;
	assign w1026 = w1791 ^ w994;
	assign w1058 = w1823 ^ w1026;
	assign w1218 = w963 ^ w48153;
	assign w1249 = w994 ^ w1218;
	assign w1281 = w1026 ^ w1249;
	assign w36926 = w36851 ^ w36825;
	assign w36815 = w36873 ^ w36846;
	assign w48088 = w36814 ^ w36815;
	assign w962 = w1727 ^ w48088;
	assign w993 = w1758 ^ w962;
	assign w1025 = w1790 ^ w993;
	assign w1057 = w1822 ^ w1025;
	assign w36699 = w1055 ^ w1057;
	assign w48092 = w36842 ^ w36813;
	assign w966 = w1731 ^ w48092;
	assign w997 = w1762 ^ w966;
	assign w1029 = w1794 ^ w997;
	assign w1061 = w1826 ^ w1029;
	assign w1221 = w966 ^ w48156;
	assign w1252 = w997 ^ w1221;
	assign w36788 = w1058 ^ w1061;
	assign w36780 = w36699 ^ w36788;
	assign w36789 = w1061 ^ w1055;
	assign w48091 = ~w36926;
	assign w965 = w1730 ^ w48091;
	assign w996 = w1761 ^ w965;
	assign w1028 = w1793 ^ w996;
	assign w1060 = w1825 ^ w1028;
	assign w36702 = w1058 ^ w1060;
	assign w484 = w1218 ^ w48217;
	assign w515 = w1249 ^ w484;
	assign w1313 = w1058 ^ w1281;
	assign w1217 = w962 ^ w48152;
	assign w1248 = w993 ^ w1217;
	assign w1280 = w1025 ^ w1248;
	assign w483 = w1217 ^ w48216;
	assign w514 = w1248 ^ w483;
	assign w1284 = w1029 ^ w1252;
	assign w1316 = w1061 ^ w1284;
	assign w36520 = w1313 ^ w1316;
	assign w36521 = w1316 ^ w1310;
	assign w546 = w1280 ^ w514;
	assign w1220 = w965 ^ w48155;
	assign w1251 = w996 ^ w1220;
	assign w1283 = w1028 ^ w1251;
	assign w1315 = w1060 ^ w1283;
	assign w36434 = w1313 ^ w1315;
	assign w486 = w1220 ^ w48219;
	assign w517 = w1251 ^ w486;
	assign w549 = w1283 ^ w517;
	assign w581 = w1315 ^ w549;
	assign w1312 = w1057 ^ w1280;
	assign w36431 = w1310 ^ w1312;
	assign w36512 = w36431 ^ w36520;
	assign w578 = w1312 ^ w546;
	assign w4903 = w576 ^ w578;
	assign w547 = w1281 ^ w515;
	assign w579 = w1313 ^ w547;
	assign w4906 = w579 ^ w581;
	assign w487 = w1221 ^ w48220;
	assign w518 = w1252 ^ w487;
	assign w550 = w1284 ^ w518;
	assign w582 = w1316 ^ w550;
	assign w4992 = w579 ^ w582;
	assign w4984 = w4903 ^ w4992;
	assign w4993 = w582 ^ w576;
	assign w44917 = w36873 ^ w36875;
	assign w36831 = w44917 ^ w36828;
	assign w36928 = w36830 ^ w36831;
	assign w48085 = ~w36928;
	assign w959 = w1724 ^ w48085;
	assign w1214 = w959 ^ w48149;
	assign w480 = w1214 ^ w48213;
	assign w990 = w1755 ^ w959;
	assign w1245 = w990 ^ w1214;
	assign w511 = w1245 ^ w480;
	assign w1022 = w1787 ^ w990;
	assign w1277 = w1022 ^ w1245;
	assign w543 = w1277 ^ w511;
	assign w1054 = w1819 ^ w1022;
	assign w36706 = w1054 ^ w1060;
	assign w1309 = w1054 ^ w1277;
	assign w36511 = w1309 ^ w36512;
	assign w36438 = w1309 ^ w1315;
	assign w575 = w1309 ^ w543;
	assign w4910 = w575 ^ w581;
	assign w36779 = w1054 ^ w36780;
	assign w4983 = w575 ^ w4984;
	assign w36818 = w36822 ^ w44917;
	assign w36821 = w36860 ^ w36818;
	assign w36925 = w36820 ^ w36821;
	assign w36817 = w36841 ^ w36818;
	assign w48087 = w36816 ^ w36817;
	assign w961 = w1726 ^ w48087;
	assign w992 = w1757 ^ w961;
	assign w1024 = w1789 ^ w992;
	assign w1056 = w1821 ^ w1024;
	assign w1216 = w961 ^ w48151;
	assign w1247 = w992 ^ w1216;
	assign w36701 = w1056 ^ w36699;
	assign w36777 = w1060 ^ w36701;
	assign w36776 = w36706 ^ w36701;
	assign w36716 = w1055 ^ w1056;
	assign w36784 = w36788 ^ w36716;
	assign w36790 = w1056 ^ w1058;
	assign w36676 = w1057 ^ w1056;
	assign w36787 = w1061 ^ w1056;
	assign w36773 = w36780 & w36784;
	assign w36705 = w36773 ^ w36702;
	assign w36767 = w36788 & w36777;
	assign w36703 = w36767 ^ w36701;
	assign w36709 = w36705 ^ w36703;
	assign w36714 = w1061 ^ w36709;
	assign w48090 = ~w36925;
	assign w964 = w1729 ^ w48090;
	assign w1219 = w964 ^ w48154;
	assign w995 = w1760 ^ w964;
	assign w1250 = w995 ^ w1219;
	assign w1027 = w1792 ^ w995;
	assign w1059 = w1824 ^ w1027;
	assign w1282 = w1027 ^ w1250;
	assign w36774 = w1059 ^ w36701;
	assign w36700 = w1059 ^ w1061;
	assign w36775 = w36700 ^ w36790;
	assign w36783 = w36700 ^ w36706;
	assign w36781 = w36716 ^ w36783;
	assign w36786 = w1059 ^ w36706;
	assign w36782 = w1055 ^ w36786;
	assign w36662 = w36702 ^ w36700;
	assign w36778 = w36699 ^ w36662;
	assign w36661 = w36702 ^ w1059;
	assign w36785 = w1054 ^ w36661;
	assign w36772 = w36781 & w36779;
	assign w36771 = w36785 & w1054;
	assign w36770 = w36789 & w36774;
	assign w36704 = w36770 ^ w36700;
	assign w36769 = w36786 & w36782;
	assign w36768 = w36783 & w36776;
	assign w36766 = w36790 & w36775;
	assign w36723 = w36766 ^ w36772;
	assign w36764 = w36723 ^ w36714;
	assign w36675 = w36766 ^ w36767;
	assign w36722 = w36675 ^ w36676;
	assign w36721 = w36722 ^ w36704;
	assign w36763 = w36769 ^ w36721;
	assign w36765 = w36787 & w36778;
	assign w36760 = w36764 & w36763;
	assign w485 = w1219 ^ w48218;
	assign w516 = w1250 ^ w485;
	assign w548 = w1282 ^ w516;
	assign w482 = w1216 ^ w48215;
	assign w513 = w1247 ^ w482;
	assign w1314 = w1059 ^ w1282;
	assign w36432 = w1314 ^ w1316;
	assign w36515 = w36432 ^ w36438;
	assign w36518 = w1314 ^ w36438;
	assign w36514 = w1310 ^ w36518;
	assign w36394 = w36434 ^ w36432;
	assign w36510 = w36431 ^ w36394;
	assign w36393 = w36434 ^ w1314;
	assign w36517 = w1309 ^ w36393;
	assign w36503 = w36517 & w1309;
	assign w36501 = w36518 & w36514;
	assign w580 = w1314 ^ w548;
	assign w4904 = w580 ^ w582;
	assign w4990 = w580 ^ w4910;
	assign w4987 = w4904 ^ w4910;
	assign w4986 = w576 ^ w4990;
	assign w4866 = w4906 ^ w4904;
	assign w4982 = w4903 ^ w4866;
	assign w4865 = w4906 ^ w580;
	assign w4973 = w4990 & w4986;
	assign w1279 = w1024 ^ w1247;
	assign w1311 = w1056 ^ w1279;
	assign w36433 = w1311 ^ w36431;
	assign w36509 = w1315 ^ w36433;
	assign w36506 = w1314 ^ w36433;
	assign w36508 = w36438 ^ w36433;
	assign w36448 = w1310 ^ w1311;
	assign w36513 = w36448 ^ w36515;
	assign w36516 = w36520 ^ w36448;
	assign w36522 = w1311 ^ w1313;
	assign w36507 = w36432 ^ w36522;
	assign w36408 = w1312 ^ w1311;
	assign w36519 = w1316 ^ w1311;
	assign w36505 = w36512 & w36516;
	assign w36437 = w36505 ^ w36434;
	assign w36504 = w36513 & w36511;
	assign w36502 = w36521 & w36506;
	assign w36436 = w36502 ^ w36432;
	assign w36500 = w36515 & w36508;
	assign w36499 = w36520 & w36509;
	assign w36435 = w36499 ^ w36433;
	assign w36441 = w36437 ^ w36435;
	assign w36446 = w1316 ^ w36441;
	assign w36498 = w36522 & w36507;
	assign w36455 = w36498 ^ w36504;
	assign w36496 = w36455 ^ w36446;
	assign w36407 = w36498 ^ w36499;
	assign w36454 = w36407 ^ w36408;
	assign w36453 = w36454 ^ w36436;
	assign w36495 = w36501 ^ w36453;
	assign w36497 = w36519 & w36510;
	assign w36492 = w36496 & w36495;
	assign w545 = w1279 ^ w513;
	assign w577 = w1311 ^ w545;
	assign w4994 = w577 ^ w579;
	assign w4979 = w4904 ^ w4994;
	assign w4920 = w576 ^ w577;
	assign w4985 = w4920 ^ w4987;
	assign w4905 = w577 ^ w4903;
	assign w4981 = w581 ^ w4905;
	assign w4980 = w4910 ^ w4905;
	assign w4978 = w580 ^ w4905;
	assign w4974 = w4993 & w4978;
	assign w4908 = w4974 ^ w4904;
	assign w4880 = w578 ^ w577;
	assign w4976 = w4985 & w4983;
	assign w4988 = w4992 ^ w4920;
	assign w4977 = w4984 & w4988;
	assign w4909 = w4977 ^ w4906;
	assign w4991 = w582 ^ w577;
	assign w4972 = w4987 & w4980;
	assign w4971 = w4992 & w4981;
	assign w4907 = w4971 ^ w4905;
	assign w4913 = w4909 ^ w4907;
	assign w4918 = w582 ^ w4913;
	assign w4970 = w4994 & w4979;
	assign w4879 = w4970 ^ w4971;
	assign w4926 = w4879 ^ w4880;
	assign w4925 = w4926 ^ w4908;
	assign w4967 = w4973 ^ w4925;
	assign w4969 = w4991 & w4982;
	assign w4927 = w4970 ^ w4976;
	assign w4968 = w4927 ^ w4918;
	assign w4964 = w4968 & w4967;
	assign w43737 = w4969 ^ w4972;
	assign w4922 = w4970 ^ w43737;
	assign w4878 = w4973 ^ w4922;
	assign w4960 = w576 ^ w4878;
	assign w4882 = w4908 ^ w43737;
	assign w4966 = w4882 ^ w4907;
	assign w4963 = w4964 ^ w4966;
	assign w4989 = w575 ^ w4865;
	assign w4975 = w4989 & w575;
	assign w43736 = w4969 ^ w4975;
	assign w4919 = w43736 ^ w4904;
	assign w4965 = w4927 ^ w4919;
	assign w4962 = w4965 & w4963;
	assign w4870 = w4962 ^ w4918;
	assign w4873 = w4962 ^ w4974;
	assign w4869 = w4873 ^ w4909;
	assign w4868 = w580 ^ w4869;
	assign w4881 = w4913 ^ w43736;
	assign w4924 = w580 ^ w4881;
	assign w4959 = w4964 ^ w4924;
	assign w4961 = w4962 ^ w4924;
	assign w4958 = w4959 & w4960;
	assign w4956 = w4964 ^ w4958;
	assign w4957 = w4958 ^ w4966;
	assign w4877 = w4958 ^ w4922;
	assign w4876 = w4958 ^ w4975;
	assign w4871 = w4876 ^ w4972;
	assign w4955 = w4966 & w4956;
	assign w4953 = w4955 ^ w4963;
	assign w4952 = w4961 & w4953;
	assign w4917 = w4952 ^ w4927;
	assign w4951 = w4917 ^ w4919;
	assign w4948 = w4917 ^ w4870;
	assign w4942 = w4948 & w4978;
	assign w4931 = w4961 & w4987;
	assign w4943 = w4957 & w575;
	assign w4875 = w4952 ^ w4976;
	assign w4941 = w4951 & w4990;
	assign w4940 = w4961 & w4980;
	assign w4884 = w4940 ^ w4941;
	assign w4934 = w4957 & w4989;
	assign w4933 = w4948 & w4993;
	assign w4900 = w4942 ^ w4933;
	assign w4932 = w4951 & w4986;
	assign w4902 = w4940 ^ w4932;
	assign w43738 = w4941 ^ w4942;
	assign w43740 = w4955 ^ w4973;
	assign w4914 = w576 ^ w43740;
	assign w4867 = w4914 ^ w4875;
	assign w4946 = w4867 ^ w4868;
	assign w4874 = w4904 ^ w4867;
	assign w4929 = w4946 & w4994;
	assign w4950 = w4871 ^ w4874;
	assign w4938 = w4946 & w4979;
	assign w4923 = w4938 ^ w43738;
	assign w4899 = w4938 ^ w4941;
	assign w4896 = ~w4899;
	assign w4937 = w4950 & w4982;
	assign w4954 = w4914 ^ w4877;
	assign w4944 = w4954 & w4983;
	assign w4935 = w4954 & w4985;
	assign w4889 = w4934 ^ w4923;
	assign w4886 = ~w4889;
	assign w4928 = w4950 & w4991;
	assign w4947 = w43740 ^ w4925;
	assign w4945 = w4947 & w4984;
	assign w4936 = w4947 & w4988;
	assign w43739 = w4943 ^ w4945;
	assign w4915 = w4933 ^ w4937;
	assign w4893 = ~w4915;
	assign w4892 = w4893 ^ w4931;
	assign w4888 = w4892 ^ w43739;
	assign w4872 = w582 ^ w4869;
	assign w4949 = w4871 ^ w4872;
	assign w4939 = w4949 & w4981;
	assign w4895 = w4938 ^ w4939;
	assign w4883 = w4939 ^ w4923;
	assign w4894 = w4939 ^ w4928;
	assign w4890 = ~w4894;
	assign w4930 = w4949 & w4992;
	assign w4891 = w4930 ^ w4888;
	assign w4995 = w4890 ^ w4891;
	assign w48250 = ~w4995;
	assign w43520 = w4929 ^ w4930;
	assign w4898 = w4902 ^ w43520;
	assign w4901 = w43739 ^ w4898;
	assign w4897 = w4893 ^ w4898;
	assign w4998 = w4900 ^ w4901;
	assign w4997 = w4896 ^ w4897;
	assign w48246 = ~w4997;
	assign w48245 = ~w4998;
	assign w4911 = w4935 ^ w43520;
	assign w4887 = w4911 ^ w4888;
	assign w48247 = w4886 ^ w4887;
	assign w4912 = w4936 ^ w4911;
	assign w4916 = w4944 ^ w4912;
	assign w4921 = w4945 ^ w4916;
	assign w48249 = w43738 ^ w4921;
	assign w4996 = w4921 ^ w4895;
	assign w48251 = ~w4996;
	assign w4885 = w4943 ^ w4916;
	assign w48248 = w4884 ^ w4885;
	assign w48252 = w4912 ^ w4883;
	assign w44897 = w36497 ^ w36503;
	assign w36447 = w44897 ^ w36432;
	assign w36493 = w36455 ^ w36447;
	assign w36409 = w36441 ^ w44897;
	assign w36452 = w1314 ^ w36409;
	assign w36487 = w36492 ^ w36452;
	assign w44898 = w36497 ^ w36500;
	assign w36450 = w36498 ^ w44898;
	assign w36406 = w36501 ^ w36450;
	assign w36488 = w1310 ^ w36406;
	assign w36486 = w36487 & w36488;
	assign w36484 = w36492 ^ w36486;
	assign w36405 = w36486 ^ w36450;
	assign w36404 = w36486 ^ w36503;
	assign w36399 = w36404 ^ w36500;
	assign w36410 = w36436 ^ w44898;
	assign w36494 = w36410 ^ w36435;
	assign w36485 = w36486 ^ w36494;
	assign w36491 = w36492 ^ w36494;
	assign w36490 = w36493 & w36491;
	assign w36489 = w36490 ^ w36452;
	assign w36401 = w36490 ^ w36502;
	assign w36397 = w36401 ^ w36437;
	assign w36400 = w1316 ^ w36397;
	assign w36477 = w36399 ^ w36400;
	assign w36398 = w36490 ^ w36446;
	assign w36396 = w1314 ^ w36397;
	assign w36483 = w36494 & w36484;
	assign w36481 = w36483 ^ w36491;
	assign w36480 = w36489 & w36481;
	assign w36445 = w36480 ^ w36455;
	assign w36479 = w36445 ^ w36447;
	assign w36403 = w36480 ^ w36504;
	assign w36476 = w36445 ^ w36398;
	assign w36471 = w36485 & w1309;
	assign w36470 = w36476 & w36506;
	assign w36469 = w36479 & w36518;
	assign w36468 = w36489 & w36508;
	assign w36412 = w36468 ^ w36469;
	assign w36467 = w36477 & w36509;
	assign w36462 = w36485 & w36517;
	assign w36461 = w36476 & w36521;
	assign w36428 = w36470 ^ w36461;
	assign w36460 = w36479 & w36514;
	assign w36430 = w36468 ^ w36460;
	assign w36459 = w36489 & w36515;
	assign w36458 = w36477 & w36520;
	assign w44899 = w36469 ^ w36470;
	assign w44901 = w36483 ^ w36501;
	assign w36442 = w1310 ^ w44901;
	assign w36395 = w36442 ^ w36403;
	assign w36402 = w36432 ^ w36395;
	assign w36478 = w36399 ^ w36402;
	assign w36474 = w36395 ^ w36396;
	assign w36466 = w36474 & w36507;
	assign w36427 = w36466 ^ w36469;
	assign w36424 = ~w36427;
	assign w36423 = w36466 ^ w36467;
	assign w36465 = w36478 & w36510;
	assign w36443 = w36461 ^ w36465;
	assign w36421 = ~w36443;
	assign w36420 = w36421 ^ w36459;
	assign w36457 = w36474 & w36522;
	assign w36456 = w36478 & w36519;
	assign w36422 = w36467 ^ w36456;
	assign w36418 = ~w36422;
	assign w43600 = w36457 ^ w36458;
	assign w36426 = w36430 ^ w43600;
	assign w36425 = w36421 ^ w36426;
	assign w36525 = w36424 ^ w36425;
	assign w48182 = ~w36525;
	assign w36482 = w36442 ^ w36405;
	assign w36472 = w36482 & w36511;
	assign w36463 = w36482 & w36513;
	assign w36439 = w36463 ^ w43600;
	assign w36451 = w36466 ^ w44899;
	assign w36417 = w36462 ^ w36451;
	assign w36414 = ~w36417;
	assign w36411 = w36467 ^ w36451;
	assign w36475 = w44901 ^ w36453;
	assign w36473 = w36475 & w36512;
	assign w36464 = w36475 & w36516;
	assign w36440 = w36464 ^ w36439;
	assign w36444 = w36472 ^ w36440;
	assign w36449 = w36473 ^ w36444;
	assign w48185 = w44899 ^ w36449;
	assign w36524 = w36449 ^ w36423;
	assign w36413 = w36471 ^ w36444;
	assign w48184 = w36412 ^ w36413;
	assign w48188 = w36440 ^ w36411;
	assign w48187 = ~w36524;
	assign w44900 = w36471 ^ w36473;
	assign w36429 = w44900 ^ w36426;
	assign w36526 = w36428 ^ w36429;
	assign w48181 = ~w36526;
	assign w36416 = w36420 ^ w44900;
	assign w36419 = w36458 ^ w36416;
	assign w36523 = w36418 ^ w36419;
	assign w36415 = w36439 ^ w36416;
	assign w48183 = w36414 ^ w36415;
	assign w48186 = ~w36523;
	assign w44908 = w36765 ^ w36768;
	assign w36678 = w36704 ^ w44908;
	assign w36762 = w36678 ^ w36703;
	assign w36759 = w36760 ^ w36762;
	assign w36718 = w36766 ^ w44908;
	assign w36674 = w36769 ^ w36718;
	assign w36756 = w1055 ^ w36674;
	assign w44911 = w36765 ^ w36771;
	assign w36677 = w36709 ^ w44911;
	assign w36720 = w1059 ^ w36677;
	assign w36755 = w36760 ^ w36720;
	assign w36754 = w36755 & w36756;
	assign w36753 = w36754 ^ w36762;
	assign w36752 = w36760 ^ w36754;
	assign w36673 = w36754 ^ w36718;
	assign w36672 = w36754 ^ w36771;
	assign w36667 = w36672 ^ w36768;
	assign w36751 = w36762 & w36752;
	assign w36749 = w36751 ^ w36759;
	assign w36739 = w36753 & w1054;
	assign w36730 = w36753 & w36785;
	assign w44910 = w36751 ^ w36769;
	assign w36743 = w44910 ^ w36721;
	assign w36741 = w36743 & w36780;
	assign w36732 = w36743 & w36784;
	assign w36710 = w1055 ^ w44910;
	assign w36750 = w36710 ^ w36673;
	assign w36740 = w36750 & w36779;
	assign w36731 = w36750 & w36781;
	assign w36715 = w44911 ^ w36700;
	assign w36761 = w36723 ^ w36715;
	assign w36758 = w36761 & w36759;
	assign w36757 = w36758 ^ w36720;
	assign w36669 = w36758 ^ w36770;
	assign w36665 = w36669 ^ w36705;
	assign w36668 = w1061 ^ w36665;
	assign w36745 = w36667 ^ w36668;
	assign w36666 = w36758 ^ w36714;
	assign w36664 = w1059 ^ w36665;
	assign w36748 = w36757 & w36749;
	assign w36713 = w36748 ^ w36723;
	assign w36747 = w36713 ^ w36715;
	assign w36671 = w36748 ^ w36772;
	assign w36663 = w36710 ^ w36671;
	assign w36670 = w36700 ^ w36663;
	assign w36746 = w36667 ^ w36670;
	assign w36744 = w36713 ^ w36666;
	assign w36742 = w36663 ^ w36664;
	assign w36738 = w36744 & w36774;
	assign w36737 = w36747 & w36786;
	assign w36736 = w36757 & w36776;
	assign w36680 = w36736 ^ w36737;
	assign w36735 = w36745 & w36777;
	assign w36734 = w36742 & w36775;
	assign w36695 = w36734 ^ w36737;
	assign w36692 = ~w36695;
	assign w36691 = w36734 ^ w36735;
	assign w36733 = w36746 & w36778;
	assign w36729 = w36744 & w36789;
	assign w36711 = w36729 ^ w36733;
	assign w36696 = w36738 ^ w36729;
	assign w36689 = ~w36711;
	assign w36728 = w36747 & w36782;
	assign w36698 = w36736 ^ w36728;
	assign w36727 = w36757 & w36783;
	assign w36688 = w36689 ^ w36727;
	assign w36726 = w36745 & w36788;
	assign w36725 = w36742 & w36790;
	assign w36724 = w36746 & w36787;
	assign w36690 = w36735 ^ w36724;
	assign w36686 = ~w36690;
	assign w44909 = w36725 ^ w36726;
	assign w36694 = w36698 ^ w44909;
	assign w36693 = w36689 ^ w36694;
	assign w36793 = w36692 ^ w36693;
	assign w48118 = ~w36793;
	assign w1087 = w1852 ^ w48118;
	assign w1119 = w864 ^ w1087;
	assign w1342 = w1087 ^ w48182;
	assign w608 = w1342 ^ w48246;
	assign w385 = w1119 ^ w1342;
	assign w1151 = w896 ^ w1119;
	assign w417 = w1151 ^ w385;
	assign w1183 = w928 ^ w1151;
	assign w449 = w1183 ^ w417;
	assign w640 = w385 ^ w608;
	assign w672 = w417 ^ w640;
	assign w704 = w449 ^ w672;
	assign w36707 = w36731 ^ w44909;
	assign w36708 = w36732 ^ w36707;
	assign w36712 = w36740 ^ w36708;
	assign w36717 = w36741 ^ w36712;
	assign w36792 = w36717 ^ w36691;
	assign w36681 = w36739 ^ w36712;
	assign w48120 = w36680 ^ w36681;
	assign w1089 = w1854 ^ w48120;
	assign w1121 = w866 ^ w1089;
	assign w48123 = ~w36792;
	assign w1092 = w1857 ^ w48123;
	assign w1124 = w869 ^ w1092;
	assign w1347 = w1092 ^ w48187;
	assign w1344 = w1089 ^ w48184;
	assign w610 = w1344 ^ w48248;
	assign w613 = w1347 ^ w48251;
	assign w387 = w1121 ^ w1344;
	assign w390 = w1124 ^ w1347;
	assign w645 = w390 ^ w613;
	assign w1156 = w901 ^ w1124;
	assign w422 = w1156 ^ w390;
	assign w677 = w422 ^ w645;
	assign w1188 = w933 ^ w1156;
	assign w454 = w1188 ^ w422;
	assign w709 = w454 ^ w677;
	assign w642 = w387 ^ w610;
	assign w1153 = w898 ^ w1121;
	assign w419 = w1153 ^ w387;
	assign w674 = w419 ^ w642;
	assign w1185 = w930 ^ w1153;
	assign w451 = w1185 ^ w419;
	assign w22361 = w449 ^ w451;
	assign w22629 = w1183 ^ w1185;
	assign w706 = w451 ^ w674;
	assign w22093 = w704 ^ w706;
	assign w44912 = w36737 ^ w36738;
	assign w48121 = w44912 ^ w36717;
	assign w1090 = w1855 ^ w48121;
	assign w1345 = w1090 ^ w48185;
	assign w611 = w1345 ^ w48249;
	assign w1122 = w867 ^ w1090;
	assign w388 = w1122 ^ w1345;
	assign w643 = w388 ^ w611;
	assign w1154 = w899 ^ w1122;
	assign w420 = w1154 ^ w388;
	assign w1186 = w931 ^ w1154;
	assign w22632 = w1186 ^ w1188;
	assign w452 = w1186 ^ w420;
	assign w22364 = w452 ^ w454;
	assign w675 = w420 ^ w643;
	assign w707 = w452 ^ w675;
	assign w22096 = w707 ^ w709;
	assign w36719 = w36734 ^ w44912;
	assign w36685 = w36730 ^ w36719;
	assign w36682 = ~w36685;
	assign w36679 = w36735 ^ w36719;
	assign w48124 = w36708 ^ w36679;
	assign w1093 = w1858 ^ w48124;
	assign w1125 = w870 ^ w1093;
	assign w1348 = w1093 ^ w48188;
	assign w391 = w1125 ^ w1348;
	assign w614 = w1348 ^ w48252;
	assign w646 = w391 ^ w614;
	assign w1157 = w902 ^ w1125;
	assign w423 = w1157 ^ w391;
	assign w678 = w423 ^ w646;
	assign w1189 = w934 ^ w1157;
	assign w22718 = w1186 ^ w1189;
	assign w22710 = w22629 ^ w22718;
	assign w22719 = w1189 ^ w1183;
	assign w455 = w1189 ^ w423;
	assign w22450 = w452 ^ w455;
	assign w22442 = w22361 ^ w22450;
	assign w22451 = w455 ^ w449;
	assign w710 = w455 ^ w678;
	assign w22182 = w707 ^ w710;
	assign w22174 = w22093 ^ w22182;
	assign w22183 = w710 ^ w704;
	assign w44913 = w36739 ^ w36741;
	assign w36697 = w44913 ^ w36694;
	assign w36794 = w36696 ^ w36697;
	assign w48117 = ~w36794;
	assign w1086 = w1851 ^ w48117;
	assign w1341 = w1086 ^ w48181;
	assign w607 = w1341 ^ w48245;
	assign w1118 = w863 ^ w1086;
	assign w1150 = w895 ^ w1118;
	assign w1182 = w927 ^ w1150;
	assign w22709 = w1182 ^ w22710;
	assign w22636 = w1182 ^ w1188;
	assign w384 = w1118 ^ w1341;
	assign w416 = w1150 ^ w384;
	assign w448 = w1182 ^ w416;
	assign w22368 = w448 ^ w454;
	assign w22441 = w448 ^ w22442;
	assign w639 = w384 ^ w607;
	assign w671 = w416 ^ w639;
	assign w703 = w448 ^ w671;
	assign w22100 = w703 ^ w709;
	assign w22173 = w703 ^ w22174;
	assign w36684 = w36688 ^ w44913;
	assign w36687 = w36726 ^ w36684;
	assign w36791 = w36686 ^ w36687;
	assign w36683 = w36707 ^ w36684;
	assign w48119 = w36682 ^ w36683;
	assign w1088 = w1853 ^ w48119;
	assign w1120 = w865 ^ w1088;
	assign w48122 = ~w36791;
	assign w1091 = w1856 ^ w48122;
	assign w1123 = w868 ^ w1091;
	assign w1343 = w1088 ^ w48183;
	assign w386 = w1120 ^ w1343;
	assign w609 = w1343 ^ w48247;
	assign w1346 = w1091 ^ w48186;
	assign w389 = w1123 ^ w1346;
	assign w612 = w1346 ^ w48250;
	assign w644 = w389 ^ w612;
	assign w1155 = w900 ^ w1123;
	assign w421 = w1155 ^ w389;
	assign w676 = w421 ^ w644;
	assign w1187 = w932 ^ w1155;
	assign w453 = w1187 ^ w421;
	assign w22362 = w453 ^ w455;
	assign w22445 = w22362 ^ w22368;
	assign w22448 = w453 ^ w22368;
	assign w22444 = w449 ^ w22448;
	assign w22324 = w22364 ^ w22362;
	assign w22440 = w22361 ^ w22324;
	assign w22323 = w22364 ^ w453;
	assign w22447 = w448 ^ w22323;
	assign w22433 = w22447 & w448;
	assign w22431 = w22448 & w22444;
	assign w22630 = w1187 ^ w1189;
	assign w22713 = w22630 ^ w22636;
	assign w22716 = w1187 ^ w22636;
	assign w22712 = w1183 ^ w22716;
	assign w22592 = w22632 ^ w22630;
	assign w22708 = w22629 ^ w22592;
	assign w22591 = w22632 ^ w1187;
	assign w22715 = w1182 ^ w22591;
	assign w22701 = w22715 & w1182;
	assign w22699 = w22716 & w22712;
	assign w708 = w453 ^ w676;
	assign w22094 = w708 ^ w710;
	assign w22177 = w22094 ^ w22100;
	assign w22180 = w708 ^ w22100;
	assign w22176 = w704 ^ w22180;
	assign w22056 = w22096 ^ w22094;
	assign w22172 = w22093 ^ w22056;
	assign w22055 = w22096 ^ w708;
	assign w22179 = w703 ^ w22055;
	assign w22165 = w703 & w22179;
	assign w22163 = w22180 & w22176;
	assign w641 = w386 ^ w609;
	assign w1152 = w897 ^ w1120;
	assign w418 = w1152 ^ w386;
	assign w673 = w418 ^ w641;
	assign w1184 = w929 ^ w1152;
	assign w22631 = w1184 ^ w22629;
	assign w22707 = w1188 ^ w22631;
	assign w22704 = w1187 ^ w22631;
	assign w22706 = w22636 ^ w22631;
	assign w22646 = w1183 ^ w1184;
	assign w22711 = w22646 ^ w22713;
	assign w22714 = w22718 ^ w22646;
	assign w22720 = w1184 ^ w1186;
	assign w22705 = w22630 ^ w22720;
	assign w22606 = w1185 ^ w1184;
	assign w22717 = w1189 ^ w1184;
	assign w22703 = w22710 & w22714;
	assign w22635 = w22703 ^ w22632;
	assign w22702 = w22711 & w22709;
	assign w22700 = w22719 & w22704;
	assign w22634 = w22700 ^ w22630;
	assign w22698 = w22713 & w22706;
	assign w22697 = w22718 & w22707;
	assign w22633 = w22697 ^ w22631;
	assign w22639 = w22635 ^ w22633;
	assign w22644 = w1189 ^ w22639;
	assign w22696 = w22720 & w22705;
	assign w22653 = w22696 ^ w22702;
	assign w22694 = w22653 ^ w22644;
	assign w22605 = w22696 ^ w22697;
	assign w22652 = w22605 ^ w22606;
	assign w22651 = w22652 ^ w22634;
	assign w22693 = w22699 ^ w22651;
	assign w22695 = w22717 & w22708;
	assign w22690 = w22694 & w22693;
	assign w450 = w1184 ^ w418;
	assign w22363 = w450 ^ w22361;
	assign w22439 = w454 ^ w22363;
	assign w22436 = w453 ^ w22363;
	assign w22438 = w22368 ^ w22363;
	assign w22378 = w449 ^ w450;
	assign w22443 = w22378 ^ w22445;
	assign w22446 = w22450 ^ w22378;
	assign w22452 = w450 ^ w452;
	assign w22437 = w22362 ^ w22452;
	assign w22338 = w451 ^ w450;
	assign w22449 = w455 ^ w450;
	assign w22435 = w22442 & w22446;
	assign w22367 = w22435 ^ w22364;
	assign w22434 = w22443 & w22441;
	assign w22432 = w22451 & w22436;
	assign w22366 = w22432 ^ w22362;
	assign w22430 = w22445 & w22438;
	assign w22429 = w22450 & w22439;
	assign w22365 = w22429 ^ w22363;
	assign w22371 = w22367 ^ w22365;
	assign w22376 = w455 ^ w22371;
	assign w22428 = w22452 & w22437;
	assign w22385 = w22428 ^ w22434;
	assign w22426 = w22385 ^ w22376;
	assign w22337 = w22428 ^ w22429;
	assign w22384 = w22337 ^ w22338;
	assign w22383 = w22384 ^ w22366;
	assign w22425 = w22431 ^ w22383;
	assign w22427 = w22449 & w22440;
	assign w22422 = w22426 & w22425;
	assign w705 = w450 ^ w673;
	assign w22095 = w705 ^ w22093;
	assign w22171 = w709 ^ w22095;
	assign w22168 = w708 ^ w22095;
	assign w22170 = w22100 ^ w22095;
	assign w22110 = w704 ^ w705;
	assign w22175 = w22110 ^ w22177;
	assign w22178 = w22182 ^ w22110;
	assign w22184 = w705 ^ w707;
	assign w22169 = w22094 ^ w22184;
	assign w22070 = w706 ^ w705;
	assign w22181 = w710 ^ w705;
	assign w22167 = w22174 & w22178;
	assign w22099 = w22167 ^ w22096;
	assign w22166 = w22175 & w22173;
	assign w22164 = w22183 & w22168;
	assign w22098 = w22164 ^ w22094;
	assign w22162 = w22177 & w22170;
	assign w22161 = w22182 & w22171;
	assign w22097 = w22161 ^ w22095;
	assign w22103 = w22099 ^ w22097;
	assign w22108 = w710 ^ w22103;
	assign w22160 = w22184 & w22169;
	assign w22117 = w22160 ^ w22166;
	assign w22158 = w22117 ^ w22108;
	assign w22069 = w22160 ^ w22161;
	assign w22116 = w22069 ^ w22070;
	assign w22115 = w22116 ^ w22098;
	assign w22157 = w22163 ^ w22115;
	assign w22159 = w22181 & w22172;
	assign w22154 = w22158 & w22157;
	assign w44295 = w22159 ^ w22165;
	assign w22109 = w44295 ^ w22094;
	assign w22155 = w22117 ^ w22109;
	assign w22071 = w22103 ^ w44295;
	assign w22114 = w708 ^ w22071;
	assign w22149 = w22154 ^ w22114;
	assign w44296 = w22159 ^ w22162;
	assign w22112 = w22160 ^ w44296;
	assign w22068 = w22163 ^ w22112;
	assign w22150 = w704 ^ w22068;
	assign w22148 = w22149 & w22150;
	assign w22146 = w22154 ^ w22148;
	assign w22067 = w22148 ^ w22112;
	assign w22066 = w22148 ^ w22165;
	assign w22061 = w22066 ^ w22162;
	assign w22072 = w22098 ^ w44296;
	assign w22156 = w22072 ^ w22097;
	assign w22147 = w22148 ^ w22156;
	assign w22153 = w22154 ^ w22156;
	assign w22152 = w22155 & w22153;
	assign w22151 = w22152 ^ w22114;
	assign w22063 = w22152 ^ w22164;
	assign w22059 = w22063 ^ w22099;
	assign w22062 = w710 ^ w22059;
	assign w22139 = w22061 ^ w22062;
	assign w22060 = w22152 ^ w22108;
	assign w22058 = w708 ^ w22059;
	assign w22145 = w22156 & w22146;
	assign w22143 = w22145 ^ w22153;
	assign w22142 = w22151 & w22143;
	assign w22107 = w22142 ^ w22117;
	assign w22141 = w22107 ^ w22109;
	assign w22065 = w22142 ^ w22166;
	assign w22138 = w22107 ^ w22060;
	assign w22133 = w22147 & w703;
	assign w22132 = w22138 & w22168;
	assign w22131 = w22141 & w22180;
	assign w22130 = w22151 & w22170;
	assign w22074 = w22130 ^ w22131;
	assign w22129 = w22139 & w22171;
	assign w22124 = w22147 & w22179;
	assign w22123 = w22138 & w22183;
	assign w22090 = w22132 ^ w22123;
	assign w22122 = w22141 & w22176;
	assign w22092 = w22130 ^ w22122;
	assign w22121 = w22151 & w22177;
	assign w22120 = w22139 & w22182;
	assign w44297 = w22131 ^ w22132;
	assign w44299 = w22145 ^ w22163;
	assign w22104 = w704 ^ w44299;
	assign w22144 = w22104 ^ w22067;
	assign w22057 = w22104 ^ w22065;
	assign w22064 = w22094 ^ w22057;
	assign w22140 = w22061 ^ w22064;
	assign w22136 = w22057 ^ w22058;
	assign w22134 = w22144 & w22173;
	assign w22128 = w22136 & w22169;
	assign w22089 = w22128 ^ w22131;
	assign w22086 = ~w22089;
	assign w22085 = w22128 ^ w22129;
	assign w22127 = w22140 & w22172;
	assign w22125 = w22144 & w22175;
	assign w22105 = w22123 ^ w22127;
	assign w22083 = ~w22105;
	assign w22082 = w22083 ^ w22121;
	assign w22119 = w22136 & w22184;
	assign w22118 = w22140 & w22181;
	assign w22084 = w22129 ^ w22118;
	assign w22080 = ~w22084;
	assign w43560 = w22119 ^ w22120;
	assign w22088 = w22092 ^ w43560;
	assign w22087 = w22083 ^ w22088;
	assign w22187 = w22086 ^ w22087;
	assign w48286 = ~w22187;
	assign w22101 = w22125 ^ w43560;
	assign w22113 = w22128 ^ w44297;
	assign w22079 = w22124 ^ w22113;
	assign w22076 = ~w22079;
	assign w22073 = w22129 ^ w22113;
	assign w22137 = w44299 ^ w22115;
	assign w22135 = w22137 & w22174;
	assign w22126 = w22137 & w22178;
	assign w22102 = w22126 ^ w22101;
	assign w22106 = w22134 ^ w22102;
	assign w22111 = w22135 ^ w22106;
	assign w48289 = w44297 ^ w22111;
	assign w22186 = w22111 ^ w22085;
	assign w22075 = w22133 ^ w22106;
	assign w48288 = w22074 ^ w22075;
	assign w48292 = w22102 ^ w22073;
	assign w48291 = ~w22186;
	assign w44298 = w22133 ^ w22135;
	assign w22091 = w44298 ^ w22088;
	assign w22188 = w22090 ^ w22091;
	assign w48285 = ~w22188;
	assign w22078 = w22082 ^ w44298;
	assign w22081 = w22120 ^ w22078;
	assign w22185 = w22080 ^ w22081;
	assign w22077 = w22101 ^ w22078;
	assign w48287 = w22076 ^ w22077;
	assign w48290 = ~w22185;
	assign w44306 = w22427 ^ w22430;
	assign w22340 = w22366 ^ w44306;
	assign w22424 = w22340 ^ w22365;
	assign w22421 = w22422 ^ w22424;
	assign w22380 = w22428 ^ w44306;
	assign w22336 = w22431 ^ w22380;
	assign w22418 = w449 ^ w22336;
	assign w44309 = w22427 ^ w22433;
	assign w22339 = w22371 ^ w44309;
	assign w22382 = w453 ^ w22339;
	assign w22417 = w22422 ^ w22382;
	assign w22416 = w22417 & w22418;
	assign w22415 = w22416 ^ w22424;
	assign w22414 = w22422 ^ w22416;
	assign w22335 = w22416 ^ w22380;
	assign w22334 = w22416 ^ w22433;
	assign w22329 = w22334 ^ w22430;
	assign w22413 = w22424 & w22414;
	assign w22411 = w22413 ^ w22421;
	assign w22401 = w22415 & w448;
	assign w22392 = w22415 & w22447;
	assign w44308 = w22413 ^ w22431;
	assign w22405 = w44308 ^ w22383;
	assign w22403 = w22405 & w22442;
	assign w22394 = w22405 & w22446;
	assign w22372 = w449 ^ w44308;
	assign w22412 = w22372 ^ w22335;
	assign w22402 = w22412 & w22441;
	assign w22393 = w22412 & w22443;
	assign w22377 = w44309 ^ w22362;
	assign w22423 = w22385 ^ w22377;
	assign w22420 = w22423 & w22421;
	assign w22419 = w22420 ^ w22382;
	assign w22331 = w22420 ^ w22432;
	assign w22327 = w22331 ^ w22367;
	assign w22330 = w455 ^ w22327;
	assign w22407 = w22329 ^ w22330;
	assign w22328 = w22420 ^ w22376;
	assign w22326 = w453 ^ w22327;
	assign w22410 = w22419 & w22411;
	assign w22375 = w22410 ^ w22385;
	assign w22409 = w22375 ^ w22377;
	assign w22333 = w22410 ^ w22434;
	assign w22325 = w22372 ^ w22333;
	assign w22332 = w22362 ^ w22325;
	assign w22408 = w22329 ^ w22332;
	assign w22406 = w22375 ^ w22328;
	assign w22404 = w22325 ^ w22326;
	assign w22400 = w22406 & w22436;
	assign w22399 = w22409 & w22448;
	assign w22398 = w22419 & w22438;
	assign w22342 = w22398 ^ w22399;
	assign w22397 = w22407 & w22439;
	assign w22396 = w22404 & w22437;
	assign w22357 = w22396 ^ w22399;
	assign w22354 = ~w22357;
	assign w22353 = w22396 ^ w22397;
	assign w22395 = w22408 & w22440;
	assign w22391 = w22406 & w22451;
	assign w22373 = w22391 ^ w22395;
	assign w22358 = w22400 ^ w22391;
	assign w22351 = ~w22373;
	assign w22390 = w22409 & w22444;
	assign w22360 = w22398 ^ w22390;
	assign w22389 = w22419 & w22445;
	assign w22350 = w22351 ^ w22389;
	assign w22388 = w22407 & w22450;
	assign w22387 = w22404 & w22452;
	assign w22386 = w22408 & w22449;
	assign w22352 = w22397 ^ w22386;
	assign w22348 = ~w22352;
	assign w44307 = w22387 ^ w22388;
	assign w22369 = w22393 ^ w44307;
	assign w22370 = w22394 ^ w22369;
	assign w22374 = w22402 ^ w22370;
	assign w22379 = w22403 ^ w22374;
	assign w22454 = w22379 ^ w22353;
	assign w22343 = w22401 ^ w22374;
	assign w48224 = w22342 ^ w22343;
	assign w48227 = ~w22454;
	assign w22356 = w22360 ^ w44307;
	assign w22355 = w22351 ^ w22356;
	assign w22455 = w22354 ^ w22355;
	assign w48222 = ~w22455;
	assign w44310 = w22399 ^ w22400;
	assign w48225 = w44310 ^ w22379;
	assign w22381 = w22396 ^ w44310;
	assign w22347 = w22392 ^ w22381;
	assign w22344 = ~w22347;
	assign w22341 = w22397 ^ w22381;
	assign w48228 = w22370 ^ w22341;
	assign w44311 = w22401 ^ w22403;
	assign w22359 = w44311 ^ w22356;
	assign w22456 = w22358 ^ w22359;
	assign w48221 = ~w22456;
	assign w22346 = w22350 ^ w44311;
	assign w22349 = w22388 ^ w22346;
	assign w22453 = w22348 ^ w22349;
	assign w22345 = w22369 ^ w22346;
	assign w48223 = w22344 ^ w22345;
	assign w48226 = ~w22453;
	assign w44317 = w22695 ^ w22701;
	assign w22607 = w22639 ^ w44317;
	assign w22650 = w1187 ^ w22607;
	assign w22685 = w22690 ^ w22650;
	assign w22645 = w44317 ^ w22630;
	assign w22691 = w22653 ^ w22645;
	assign w44318 = w22695 ^ w22698;
	assign w22648 = w22696 ^ w44318;
	assign w22604 = w22699 ^ w22648;
	assign w22686 = w1183 ^ w22604;
	assign w22684 = w22685 & w22686;
	assign w22682 = w22690 ^ w22684;
	assign w22602 = w22684 ^ w22701;
	assign w22597 = w22602 ^ w22698;
	assign w22603 = w22684 ^ w22648;
	assign w22608 = w22634 ^ w44318;
	assign w22692 = w22608 ^ w22633;
	assign w22683 = w22684 ^ w22692;
	assign w22689 = w22690 ^ w22692;
	assign w22688 = w22691 & w22689;
	assign w22687 = w22688 ^ w22650;
	assign w22599 = w22688 ^ w22700;
	assign w22595 = w22599 ^ w22635;
	assign w22598 = w1189 ^ w22595;
	assign w22675 = w22597 ^ w22598;
	assign w22596 = w22688 ^ w22644;
	assign w22594 = w1187 ^ w22595;
	assign w22681 = w22692 & w22682;
	assign w22679 = w22681 ^ w22689;
	assign w22678 = w22687 & w22679;
	assign w22643 = w22678 ^ w22653;
	assign w22677 = w22643 ^ w22645;
	assign w22601 = w22678 ^ w22702;
	assign w22674 = w22643 ^ w22596;
	assign w22669 = w22683 & w1182;
	assign w22668 = w22674 & w22704;
	assign w22667 = w22677 & w22716;
	assign w22666 = w22687 & w22706;
	assign w22610 = w22666 ^ w22667;
	assign w22665 = w22675 & w22707;
	assign w22660 = w22683 & w22715;
	assign w22659 = w22674 & w22719;
	assign w22626 = w22668 ^ w22659;
	assign w22658 = w22677 & w22712;
	assign w22628 = w22666 ^ w22658;
	assign w22657 = w22687 & w22713;
	assign w22656 = w22675 & w22718;
	assign w44320 = w22667 ^ w22668;
	assign w44322 = w22681 ^ w22699;
	assign w22673 = w44322 ^ w22651;
	assign w22662 = w22673 & w22714;
	assign w22671 = w22673 & w22710;
	assign w44321 = w22669 ^ w22671;
	assign w22640 = w1183 ^ w44322;
	assign w22680 = w22640 ^ w22603;
	assign w22593 = w22640 ^ w22601;
	assign w22600 = w22630 ^ w22593;
	assign w22676 = w22597 ^ w22600;
	assign w22672 = w22593 ^ w22594;
	assign w22670 = w22680 & w22709;
	assign w22664 = w22672 & w22705;
	assign w22649 = w22664 ^ w44320;
	assign w22625 = w22664 ^ w22667;
	assign w22622 = ~w22625;
	assign w22621 = w22664 ^ w22665;
	assign w22615 = w22660 ^ w22649;
	assign w22612 = ~w22615;
	assign w22609 = w22665 ^ w22649;
	assign w22663 = w22676 & w22708;
	assign w22641 = w22659 ^ w22663;
	assign w22619 = ~w22641;
	assign w22618 = w22619 ^ w22657;
	assign w22614 = w22618 ^ w44321;
	assign w22617 = w22656 ^ w22614;
	assign w22661 = w22680 & w22711;
	assign w22655 = w22672 & w22720;
	assign w22654 = w22676 & w22717;
	assign w22620 = w22665 ^ w22654;
	assign w22616 = ~w22620;
	assign w22721 = w22616 ^ w22617;
	assign w48162 = ~w22721;
	assign w1227 = w972 ^ w48162;
	assign w493 = w1227 ^ w48226;
	assign w748 = w493 ^ w48290;
	assign w1258 = w1003 ^ w1227;
	assign w1290 = w1035 ^ w1258;
	assign w524 = w1258 ^ w493;
	assign w556 = w1290 ^ w524;
	assign w1322 = w1067 ^ w1290;
	assign w780 = w524 ^ w748;
	assign w588 = w1322 ^ w556;
	assign w44319 = w22655 ^ w22656;
	assign w22637 = w22661 ^ w44319;
	assign w22613 = w22637 ^ w22614;
	assign w48159 = w22612 ^ w22613;
	assign w1224 = w969 ^ w48159;
	assign w1255 = w1000 ^ w1224;
	assign w1287 = w1032 ^ w1255;
	assign w490 = w1224 ^ w48223;
	assign w1319 = w1064 ^ w1287;
	assign w521 = w1255 ^ w490;
	assign w553 = w1287 ^ w521;
	assign w585 = w1319 ^ w553;
	assign w745 = w490 ^ w48287;
	assign w777 = w521 ^ w745;
	assign w22638 = w22662 ^ w22637;
	assign w48164 = w22638 ^ w22609;
	assign w1229 = w974 ^ w48164;
	assign w1260 = w1005 ^ w1229;
	assign w1292 = w1037 ^ w1260;
	assign w1324 = w1069 ^ w1292;
	assign w22583 = w1324 ^ w1319;
	assign w22496 = w1322 ^ w1324;
	assign w22642 = w22670 ^ w22638;
	assign w22611 = w22669 ^ w22642;
	assign w48160 = w22610 ^ w22611;
	assign w1225 = w970 ^ w48160;
	assign w491 = w1225 ^ w48224;
	assign w746 = w491 ^ w48288;
	assign w1256 = w1001 ^ w1225;
	assign w522 = w1256 ^ w491;
	assign w778 = w522 ^ w746;
	assign w1288 = w1033 ^ w1256;
	assign w554 = w1288 ^ w522;
	assign w810 = w554 ^ w778;
	assign w1320 = w1065 ^ w1288;
	assign w586 = w1320 ^ w554;
	assign w22204 = w586 ^ w585;
	assign w842 = w586 ^ w810;
	assign w22472 = w1320 ^ w1319;
	assign w22647 = w22671 ^ w22642;
	assign w22722 = w22647 ^ w22621;
	assign w48163 = ~w22722;
	assign w1228 = w973 ^ w48163;
	assign w494 = w1228 ^ w48227;
	assign w1259 = w1004 ^ w1228;
	assign w1291 = w1036 ^ w1259;
	assign w1323 = w1068 ^ w1291;
	assign w525 = w1259 ^ w494;
	assign w557 = w1291 ^ w525;
	assign w589 = w1323 ^ w557;
	assign w749 = w494 ^ w48291;
	assign w781 = w525 ^ w749;
	assign w813 = w557 ^ w781;
	assign w845 = w589 ^ w813;
	assign w48161 = w44320 ^ w22647;
	assign w1226 = w971 ^ w48161;
	assign w1257 = w1002 ^ w1226;
	assign w1289 = w1034 ^ w1257;
	assign w1321 = w1066 ^ w1289;
	assign w22584 = w1321 ^ w1324;
	assign w22498 = w1321 ^ w1323;
	assign w22586 = w1319 ^ w1321;
	assign w492 = w1226 ^ w48225;
	assign w523 = w1257 ^ w492;
	assign w22571 = w22496 ^ w22586;
	assign w22458 = w22498 ^ w22496;
	assign w22457 = w22498 ^ w1322;
	assign w22562 = w22586 & w22571;
	assign w555 = w1289 ^ w523;
	assign w587 = w1321 ^ w555;
	assign w22230 = w587 ^ w589;
	assign w22189 = w22230 ^ w588;
	assign w22318 = w585 ^ w587;
	assign w747 = w492 ^ w48289;
	assign w779 = w523 ^ w747;
	assign w811 = w555 ^ w779;
	assign w843 = w587 ^ w811;
	assign w22624 = w22628 ^ w44319;
	assign w22627 = w44321 ^ w22624;
	assign w22724 = w22626 ^ w22627;
	assign w22623 = w22619 ^ w22624;
	assign w22723 = w22622 ^ w22623;
	assign w48157 = ~w22724;
	assign w48158 = ~w22723;
	assign w1223 = w968 ^ w48158;
	assign w1254 = w999 ^ w1223;
	assign w1286 = w1031 ^ w1254;
	assign w489 = w1223 ^ w48222;
	assign w1222 = w967 ^ w48157;
	assign w1253 = w998 ^ w1222;
	assign w488 = w1222 ^ w48221;
	assign w743 = w488 ^ w48285;
	assign w519 = w1253 ^ w488;
	assign w775 = w519 ^ w743;
	assign w1285 = w1030 ^ w1253;
	assign w520 = w1254 ^ w489;
	assign w552 = w1286 ^ w520;
	assign w1318 = w1063 ^ w1286;
	assign w22495 = w1318 ^ w1320;
	assign w22497 = w1319 ^ w22495;
	assign w22573 = w1323 ^ w22497;
	assign w22570 = w1322 ^ w22497;
	assign w22576 = w22495 ^ w22584;
	assign w22512 = w1318 ^ w1319;
	assign w22580 = w22584 ^ w22512;
	assign w22574 = w22495 ^ w22458;
	assign w22585 = w1324 ^ w1318;
	assign w22569 = w22576 & w22580;
	assign w22501 = w22569 ^ w22498;
	assign w22566 = w22585 & w22570;
	assign w22500 = w22566 ^ w22496;
	assign w22563 = w22584 & w22573;
	assign w22499 = w22563 ^ w22497;
	assign w22505 = w22501 ^ w22499;
	assign w22510 = w1324 ^ w22505;
	assign w22471 = w22562 ^ w22563;
	assign w22518 = w22471 ^ w22472;
	assign w22517 = w22518 ^ w22500;
	assign w22561 = w22583 & w22574;
	assign w584 = w1318 ^ w552;
	assign w22227 = w584 ^ w586;
	assign w22229 = w585 ^ w22227;
	assign w22305 = w589 ^ w22229;
	assign w22302 = w588 ^ w22229;
	assign w22244 = w584 ^ w585;
	assign w1317 = w1062 ^ w1285;
	assign w22575 = w1317 ^ w22576;
	assign w22502 = w1317 ^ w1323;
	assign w22572 = w22502 ^ w22497;
	assign w22579 = w22496 ^ w22502;
	assign w22577 = w22512 ^ w22579;
	assign w22582 = w1322 ^ w22502;
	assign w22578 = w1318 ^ w22582;
	assign w22581 = w1317 ^ w22457;
	assign w22568 = w22577 & w22575;
	assign w22519 = w22562 ^ w22568;
	assign w22560 = w22519 ^ w22510;
	assign w22567 = w22581 & w1317;
	assign w22565 = w22582 & w22578;
	assign w22559 = w22565 ^ w22517;
	assign w22564 = w22579 & w22572;
	assign w22556 = w22560 & w22559;
	assign w744 = w489 ^ w48286;
	assign w551 = w1285 ^ w519;
	assign w583 = w1317 ^ w551;
	assign w22234 = w583 ^ w589;
	assign w22304 = w22234 ^ w22229;
	assign w22314 = w588 ^ w22234;
	assign w22310 = w584 ^ w22314;
	assign w22313 = w583 ^ w22189;
	assign w22299 = w22313 & w583;
	assign w22297 = w22314 & w22310;
	assign w807 = w551 ^ w775;
	assign w839 = w583 ^ w807;
	assign w44312 = w22561 ^ w22567;
	assign w22511 = w44312 ^ w22496;
	assign w22557 = w22519 ^ w22511;
	assign w22473 = w22505 ^ w44312;
	assign w22516 = w1322 ^ w22473;
	assign w22551 = w22556 ^ w22516;
	assign w44313 = w22561 ^ w22564;
	assign w22514 = w22562 ^ w44313;
	assign w22470 = w22565 ^ w22514;
	assign w22552 = w1318 ^ w22470;
	assign w22550 = w22551 & w22552;
	assign w22548 = w22556 ^ w22550;
	assign w22469 = w22550 ^ w22514;
	assign w22468 = w22550 ^ w22567;
	assign w22463 = w22468 ^ w22564;
	assign w22474 = w22500 ^ w44313;
	assign w22558 = w22474 ^ w22499;
	assign w22549 = w22550 ^ w22558;
	assign w22555 = w22556 ^ w22558;
	assign w22554 = w22557 & w22555;
	assign w22553 = w22554 ^ w22516;
	assign w22465 = w22554 ^ w22566;
	assign w22461 = w22465 ^ w22501;
	assign w22464 = w1324 ^ w22461;
	assign w22541 = w22463 ^ w22464;
	assign w22462 = w22554 ^ w22510;
	assign w22460 = w1322 ^ w22461;
	assign w22547 = w22558 & w22548;
	assign w22545 = w22547 ^ w22555;
	assign w22544 = w22553 & w22545;
	assign w22509 = w22544 ^ w22519;
	assign w22543 = w22509 ^ w22511;
	assign w22467 = w22544 ^ w22568;
	assign w22540 = w22509 ^ w22462;
	assign w22535 = w22549 & w1317;
	assign w22534 = w22540 & w22570;
	assign w22533 = w22543 & w22582;
	assign w22532 = w22553 & w22572;
	assign w22476 = w22532 ^ w22533;
	assign w22531 = w22541 & w22573;
	assign w22526 = w22549 & w22581;
	assign w22525 = w22540 & w22585;
	assign w22492 = w22534 ^ w22525;
	assign w22524 = w22543 & w22578;
	assign w22494 = w22532 ^ w22524;
	assign w22523 = w22553 & w22579;
	assign w22522 = w22541 & w22584;
	assign w44314 = w22533 ^ w22534;
	assign w44316 = w22547 ^ w22565;
	assign w22506 = w1318 ^ w44316;
	assign w22546 = w22506 ^ w22469;
	assign w22536 = w22546 & w22575;
	assign w22527 = w22546 & w22577;
	assign w22459 = w22506 ^ w22467;
	assign w22538 = w22459 ^ w22460;
	assign w22530 = w22538 & w22571;
	assign w22491 = w22530 ^ w22533;
	assign w22488 = ~w22491;
	assign w22487 = w22530 ^ w22531;
	assign w22521 = w22538 & w22586;
	assign w43561 = w22521 ^ w22522;
	assign w22503 = w22527 ^ w43561;
	assign w22490 = w22494 ^ w43561;
	assign w22466 = w22496 ^ w22459;
	assign w22515 = w22530 ^ w44314;
	assign w22481 = w22526 ^ w22515;
	assign w22478 = ~w22481;
	assign w22475 = w22531 ^ w22515;
	assign w22542 = w22463 ^ w22466;
	assign w22520 = w22542 & w22583;
	assign w22486 = w22531 ^ w22520;
	assign w22482 = ~w22486;
	assign w22529 = w22542 & w22574;
	assign w22507 = w22525 ^ w22529;
	assign w22485 = ~w22507;
	assign w22484 = w22485 ^ w22523;
	assign w22489 = w22485 ^ w22490;
	assign w22589 = w22488 ^ w22489;
	assign w48190 = ~w22589;
	assign w1350 = w1095 ^ w48190;
	assign w393 = w1127 ^ w1350;
	assign w425 = w1159 ^ w393;
	assign w457 = w1191 ^ w425;
	assign w22539 = w44316 ^ w22517;
	assign w22537 = w22539 & w22576;
	assign w22528 = w22539 & w22580;
	assign w22504 = w22528 ^ w22503;
	assign w22508 = w22536 ^ w22504;
	assign w22513 = w22537 ^ w22508;
	assign w48193 = w44314 ^ w22513;
	assign w22588 = w22513 ^ w22487;
	assign w22477 = w22535 ^ w22508;
	assign w48192 = w22476 ^ w22477;
	assign w48196 = w22504 ^ w22475;
	assign w48195 = ~w22588;
	assign w1352 = w1097 ^ w48192;
	assign w1353 = w1098 ^ w48193;
	assign w395 = w1129 ^ w1352;
	assign w427 = w1161 ^ w395;
	assign w1356 = w1101 ^ w48196;
	assign w399 = w1133 ^ w1356;
	assign w431 = w1165 ^ w399;
	assign w463 = w1197 ^ w431;
	assign w34779 = w463 ^ w457;
	assign w1355 = w1100 ^ w48195;
	assign w398 = w1132 ^ w1355;
	assign w430 = w1164 ^ w398;
	assign w462 = w1196 ^ w430;
	assign w44315 = w22535 ^ w22537;
	assign w22493 = w44315 ^ w22490;
	assign w22590 = w22492 ^ w22493;
	assign w48189 = ~w22590;
	assign w22480 = w22484 ^ w44315;
	assign w22483 = w22522 ^ w22480;
	assign w22587 = w22482 ^ w22483;
	assign w22479 = w22503 ^ w22480;
	assign w48191 = w22478 ^ w22479;
	assign w48194 = ~w22587;
	assign w1351 = w1096 ^ w48191;
	assign w394 = w1128 ^ w1351;
	assign w426 = w1160 ^ w394;
	assign w458 = w1192 ^ w426;
	assign w34706 = w457 ^ w458;
	assign w34777 = w463 ^ w458;
	assign w1354 = w1099 ^ w48194;
	assign w397 = w1131 ^ w1354;
	assign w429 = w1163 ^ w397;
	assign w461 = w1195 ^ w429;
	assign w34690 = w461 ^ w463;
	assign w1349 = w1094 ^ w48189;
	assign w392 = w1126 ^ w1349;
	assign w424 = w1158 ^ w392;
	assign w396 = w1130 ^ w1353;
	assign w428 = w1162 ^ w396;
	assign w460 = w1194 ^ w428;
	assign w34692 = w460 ^ w462;
	assign w34778 = w460 ^ w463;
	assign w34774 = w34778 ^ w34706;
	assign w34780 = w458 ^ w460;
	assign w34765 = w34690 ^ w34780;
	assign w34652 = w34692 ^ w34690;
	assign w34651 = w34692 ^ w461;
	assign w34756 = w34780 & w34765;
	assign w495 = w1229 ^ w48228;
	assign w750 = w495 ^ w48292;
	assign w526 = w1260 ^ w495;
	assign w558 = w1292 ^ w526;
	assign w590 = w1324 ^ w558;
	assign w22228 = w588 ^ w590;
	assign w22303 = w22228 ^ w22318;
	assign w22316 = w587 ^ w590;
	assign w22312 = w22316 ^ w22244;
	assign w22311 = w22228 ^ w22234;
	assign w22309 = w22244 ^ w22311;
	assign w22308 = w22227 ^ w22316;
	assign w22307 = w583 ^ w22308;
	assign w22190 = w22230 ^ w22228;
	assign w22306 = w22227 ^ w22190;
	assign w22317 = w590 ^ w584;
	assign w22315 = w590 ^ w585;
	assign w22301 = w22308 & w22312;
	assign w22233 = w22301 ^ w22230;
	assign w22300 = w22309 & w22307;
	assign w22298 = w22317 & w22302;
	assign w22232 = w22298 ^ w22228;
	assign w22296 = w22311 & w22304;
	assign w22295 = w22316 & w22305;
	assign w22231 = w22295 ^ w22229;
	assign w22237 = w22233 ^ w22231;
	assign w22242 = w590 ^ w22237;
	assign w22294 = w22318 & w22303;
	assign w22251 = w22294 ^ w22300;
	assign w22292 = w22251 ^ w22242;
	assign w22203 = w22294 ^ w22295;
	assign w22250 = w22203 ^ w22204;
	assign w22249 = w22250 ^ w22232;
	assign w22291 = w22297 ^ w22249;
	assign w22293 = w22315 & w22306;
	assign w22288 = w22292 & w22291;
	assign w782 = w526 ^ w750;
	assign w814 = w558 ^ w782;
	assign w846 = w590 ^ w814;
	assign w44300 = w22293 ^ w22299;
	assign w22205 = w22237 ^ w44300;
	assign w22248 = w588 ^ w22205;
	assign w22283 = w22288 ^ w22248;
	assign w22243 = w44300 ^ w22228;
	assign w22289 = w22251 ^ w22243;
	assign w44301 = w22293 ^ w22296;
	assign w22246 = w22294 ^ w44301;
	assign w22202 = w22297 ^ w22246;
	assign w22284 = w584 ^ w22202;
	assign w22282 = w22283 & w22284;
	assign w22280 = w22288 ^ w22282;
	assign w22201 = w22282 ^ w22246;
	assign w22200 = w22282 ^ w22299;
	assign w22195 = w22200 ^ w22296;
	assign w22206 = w22232 ^ w44301;
	assign w22290 = w22206 ^ w22231;
	assign w22281 = w22282 ^ w22290;
	assign w22287 = w22288 ^ w22290;
	assign w22286 = w22289 & w22287;
	assign w22285 = w22286 ^ w22248;
	assign w22197 = w22286 ^ w22298;
	assign w22193 = w22197 ^ w22233;
	assign w22196 = w590 ^ w22193;
	assign w22273 = w22195 ^ w22196;
	assign w22194 = w22286 ^ w22242;
	assign w22192 = w588 ^ w22193;
	assign w22279 = w22290 & w22280;
	assign w22277 = w22279 ^ w22287;
	assign w22276 = w22285 & w22277;
	assign w22241 = w22276 ^ w22251;
	assign w22275 = w22241 ^ w22243;
	assign w22199 = w22276 ^ w22300;
	assign w22272 = w22241 ^ w22194;
	assign w22267 = w22281 & w583;
	assign w22266 = w22272 & w22302;
	assign w22265 = w22275 & w22314;
	assign w22264 = w22285 & w22304;
	assign w22208 = w22264 ^ w22265;
	assign w22263 = w22273 & w22305;
	assign w22258 = w22281 & w22313;
	assign w22257 = w22272 & w22317;
	assign w22224 = w22266 ^ w22257;
	assign w22256 = w22275 & w22310;
	assign w22226 = w22264 ^ w22256;
	assign w22255 = w22285 & w22311;
	assign w22254 = w22273 & w22316;
	assign w44303 = w22265 ^ w22266;
	assign w44305 = w22279 ^ w22297;
	assign w22271 = w44305 ^ w22249;
	assign w22260 = w22271 & w22312;
	assign w22269 = w22271 & w22308;
	assign w44304 = w22267 ^ w22269;
	assign w22238 = w584 ^ w44305;
	assign w22278 = w22238 ^ w22201;
	assign w22191 = w22238 ^ w22199;
	assign w22198 = w22228 ^ w22191;
	assign w22274 = w22195 ^ w22198;
	assign w22270 = w22191 ^ w22192;
	assign w22268 = w22278 & w22307;
	assign w22262 = w22270 & w22303;
	assign w22247 = w22262 ^ w44303;
	assign w22223 = w22262 ^ w22265;
	assign w22220 = ~w22223;
	assign w22219 = w22262 ^ w22263;
	assign w22213 = w22258 ^ w22247;
	assign w22210 = ~w22213;
	assign w22207 = w22263 ^ w22247;
	assign w22261 = w22274 & w22306;
	assign w22239 = w22257 ^ w22261;
	assign w22217 = ~w22239;
	assign w22216 = w22217 ^ w22255;
	assign w22212 = w22216 ^ w44304;
	assign w22215 = w22254 ^ w22212;
	assign w22259 = w22278 & w22309;
	assign w22253 = w22270 & w22318;
	assign w22252 = w22274 & w22315;
	assign w22218 = w22263 ^ w22252;
	assign w22214 = ~w22218;
	assign w22319 = w22214 ^ w22215;
	assign w48258 = ~w22319;
	assign w620 = w1354 ^ w48258;
	assign w652 = w397 ^ w620;
	assign w684 = w429 ^ w652;
	assign w716 = w461 ^ w684;
	assign w44302 = w22253 ^ w22254;
	assign w22235 = w22259 ^ w44302;
	assign w22236 = w22260 ^ w22235;
	assign w22240 = w22268 ^ w22236;
	assign w22245 = w22269 ^ w22240;
	assign w48257 = w44303 ^ w22245;
	assign w619 = w1353 ^ w48257;
	assign w651 = w396 ^ w619;
	assign w22320 = w22245 ^ w22219;
	assign w22211 = w22235 ^ w22212;
	assign w48255 = w22210 ^ w22211;
	assign w22209 = w22267 ^ w22240;
	assign w48256 = w22208 ^ w22209;
	assign w48260 = w22236 ^ w22207;
	assign w622 = w1356 ^ w48260;
	assign w48259 = ~w22320;
	assign w617 = w1351 ^ w48255;
	assign w649 = w394 ^ w617;
	assign w683 = w428 ^ w651;
	assign w654 = w399 ^ w622;
	assign w686 = w431 ^ w654;
	assign w718 = w463 ^ w686;
	assign w715 = w460 ^ w683;
	assign w5127 = w715 ^ w718;
	assign w681 = w426 ^ w649;
	assign w713 = w458 ^ w681;
	assign w5129 = w713 ^ w715;
	assign w5126 = w718 ^ w713;
	assign w621 = w1355 ^ w48259;
	assign w653 = w398 ^ w621;
	assign w685 = w430 ^ w653;
	assign w717 = w462 ^ w685;
	assign w5040 = w715 ^ w717;
	assign w618 = w1352 ^ w48256;
	assign w650 = w395 ^ w618;
	assign w682 = w427 ^ w650;
	assign w4999 = w5040 ^ w716;
	assign w5038 = w716 ^ w718;
	assign w5000 = w5040 ^ w5038;
	assign w5114 = w5038 ^ w5129;
	assign w5105 = w5129 & w5114;
	assign w22222 = w22226 ^ w44302;
	assign w22225 = w44304 ^ w22222;
	assign w22322 = w22224 ^ w22225;
	assign w22221 = w22217 ^ w22222;
	assign w22321 = w22220 ^ w22221;
	assign w48253 = ~w22322;
	assign w48254 = ~w22321;
	assign w616 = w1350 ^ w48254;
	assign w648 = w393 ^ w616;
	assign w680 = w425 ^ w648;
	assign w712 = w457 ^ w680;
	assign w5128 = w718 ^ w712;
	assign w5054 = w712 ^ w713;
	assign w5123 = w5127 ^ w5054;
	assign w615 = w1349 ^ w48253;
	assign w647 = w392 ^ w615;
	assign w679 = w424 ^ w647;
	assign w459 = w1193 ^ w427;
	assign w34689 = w457 ^ w459;
	assign w34691 = w458 ^ w34689;
	assign w34767 = w462 ^ w34691;
	assign w34764 = w461 ^ w34691;
	assign w34770 = w34689 ^ w34778;
	assign w34666 = w459 ^ w458;
	assign w34768 = w34689 ^ w34652;
	assign w34763 = w34770 & w34774;
	assign w34695 = w34763 ^ w34692;
	assign w34760 = w34779 & w34764;
	assign w34694 = w34760 ^ w34690;
	assign w34757 = w34778 & w34767;
	assign w34693 = w34757 ^ w34691;
	assign w34699 = w34695 ^ w34693;
	assign w34704 = w463 ^ w34699;
	assign w34665 = w34756 ^ w34757;
	assign w34712 = w34665 ^ w34666;
	assign w34711 = w34712 ^ w34694;
	assign w34755 = w34777 & w34768;
	assign w714 = w459 ^ w682;
	assign w5014 = w714 ^ w713;
	assign w5037 = w712 ^ w714;
	assign w5039 = w713 ^ w5037;
	assign w5117 = w5037 ^ w5000;
	assign w5104 = w5126 & w5117;
	assign w5113 = w716 ^ w5039;
	assign w5109 = w5128 & w5113;
	assign w5042 = w5109 ^ w5038;
	assign w5119 = w5037 ^ w5127;
	assign w5112 = w5119 & w5123;
	assign w5043 = w5112 ^ w5040;
	assign w5116 = w717 ^ w5039;
	assign w5106 = w5127 & w5116;
	assign w5041 = w5106 ^ w5039;
	assign w5013 = w5105 ^ w5106;
	assign w5060 = w5013 ^ w5014;
	assign w5059 = w5060 ^ w5042;
	assign w5047 = w5043 ^ w5041;
	assign w5052 = w718 ^ w5047;
	assign w456 = w1190 ^ w424;
	assign w34769 = w456 ^ w34770;
	assign w34696 = w456 ^ w462;
	assign w34766 = w34696 ^ w34691;
	assign w34773 = w34690 ^ w34696;
	assign w34771 = w34706 ^ w34773;
	assign w34776 = w461 ^ w34696;
	assign w34772 = w457 ^ w34776;
	assign w34775 = w456 ^ w34651;
	assign w34762 = w34771 & w34769;
	assign w34713 = w34756 ^ w34762;
	assign w34754 = w34713 ^ w34704;
	assign w34761 = w34775 & w456;
	assign w34759 = w34776 & w34772;
	assign w34753 = w34759 ^ w34711;
	assign w34758 = w34773 & w34766;
	assign w34750 = w34754 & w34753;
	assign w711 = w456 ^ w679;
	assign w5124 = w711 ^ w4999;
	assign w5110 = w711 & w5124;
	assign w5044 = w711 ^ w717;
	assign w5122 = w5038 ^ w5044;
	assign w5125 = w716 ^ w5044;
	assign w5121 = w712 ^ w5125;
	assign w5108 = w5125 & w5121;
	assign w5102 = w5108 ^ w5059;
	assign w5118 = w711 ^ w5119;
	assign w5115 = w5044 ^ w5039;
	assign w5107 = w5122 & w5115;
	assign w5120 = w5054 ^ w5122;
	assign w5111 = w5120 & w5118;
	assign w5061 = w5105 ^ w5111;
	assign w5103 = w5061 ^ w5052;
	assign w5099 = w5103 & w5102;
	assign w44823 = w34755 ^ w34758;
	assign w34668 = w34694 ^ w44823;
	assign w34752 = w34668 ^ w34693;
	assign w34749 = w34750 ^ w34752;
	assign w34708 = w34756 ^ w44823;
	assign w34664 = w34759 ^ w34708;
	assign w34746 = w457 ^ w34664;
	assign w44826 = w34755 ^ w34761;
	assign w34667 = w34699 ^ w44826;
	assign w34710 = w461 ^ w34667;
	assign w34745 = w34750 ^ w34710;
	assign w34744 = w34745 & w34746;
	assign w34743 = w34744 ^ w34752;
	assign w34742 = w34750 ^ w34744;
	assign w34663 = w34744 ^ w34708;
	assign w34662 = w34744 ^ w34761;
	assign w34657 = w34662 ^ w34758;
	assign w34741 = w34752 & w34742;
	assign w34739 = w34741 ^ w34749;
	assign w34729 = w34743 & w456;
	assign w34720 = w34743 & w34775;
	assign w44825 = w34741 ^ w34759;
	assign w34733 = w44825 ^ w34711;
	assign w34731 = w34733 & w34770;
	assign w34722 = w34733 & w34774;
	assign w34700 = w457 ^ w44825;
	assign w34740 = w34700 ^ w34663;
	assign w34730 = w34740 & w34769;
	assign w34721 = w34740 & w34771;
	assign w34705 = w44826 ^ w34690;
	assign w34751 = w34713 ^ w34705;
	assign w34748 = w34751 & w34749;
	assign w34747 = w34748 ^ w34710;
	assign w34659 = w34748 ^ w34760;
	assign w34655 = w34659 ^ w34695;
	assign w34658 = w463 ^ w34655;
	assign w34735 = w34657 ^ w34658;
	assign w34656 = w34748 ^ w34704;
	assign w34654 = w461 ^ w34655;
	assign w34738 = w34747 & w34739;
	assign w34703 = w34738 ^ w34713;
	assign w34737 = w34703 ^ w34705;
	assign w34661 = w34738 ^ w34762;
	assign w34653 = w34700 ^ w34661;
	assign w34660 = w34690 ^ w34653;
	assign w34736 = w34657 ^ w34660;
	assign w34734 = w34703 ^ w34656;
	assign w34732 = w34653 ^ w34654;
	assign w34728 = w34734 & w34764;
	assign w34727 = w34737 & w34776;
	assign w34726 = w34747 & w34766;
	assign w34670 = w34726 ^ w34727;
	assign w34725 = w34735 & w34767;
	assign w34724 = w34732 & w34765;
	assign w34685 = w34724 ^ w34727;
	assign w34682 = ~w34685;
	assign w34681 = w34724 ^ w34725;
	assign w34723 = w34736 & w34768;
	assign w34719 = w34734 & w34779;
	assign w34701 = w34719 ^ w34723;
	assign w34686 = w34728 ^ w34719;
	assign w34679 = ~w34701;
	assign w34718 = w34737 & w34772;
	assign w34688 = w34726 ^ w34718;
	assign w34717 = w34747 & w34773;
	assign w34678 = w34679 ^ w34717;
	assign w34716 = w34735 & w34778;
	assign w34715 = w34732 & w34780;
	assign w34714 = w34736 & w34777;
	assign w34680 = w34725 ^ w34714;
	assign w34676 = ~w34680;
	assign w44824 = w34715 ^ w34716;
	assign w34697 = w34721 ^ w44824;
	assign w34698 = w34722 ^ w34697;
	assign w34702 = w34730 ^ w34698;
	assign w34707 = w34731 ^ w34702;
	assign w34782 = w34707 ^ w34681;
	assign w34671 = w34729 ^ w34702;
	assign w48232 = w34670 ^ w34671;
	assign w48235 = ~w34782;
	assign w502 = w1236 ^ w48235;
	assign w499 = w1233 ^ w48232;
	assign w530 = w1264 ^ w499;
	assign w562 = w1296 ^ w530;
	assign w594 = w1328 ^ w562;
	assign w533 = w1267 ^ w502;
	assign w565 = w1299 ^ w533;
	assign w597 = w1331 ^ w565;
	assign w34684 = w34688 ^ w44824;
	assign w34683 = w34679 ^ w34684;
	assign w34783 = w34682 ^ w34683;
	assign w48230 = ~w34783;
	assign w497 = w1231 ^ w48230;
	assign w528 = w1262 ^ w497;
	assign w560 = w1294 ^ w528;
	assign w592 = w1326 ^ w560;
	assign w34555 = w592 ^ w594;
	assign w44827 = w34727 ^ w34728;
	assign w48233 = w44827 ^ w34707;
	assign w500 = w1234 ^ w48233;
	assign w531 = w1265 ^ w500;
	assign w563 = w1297 ^ w531;
	assign w595 = w1329 ^ w563;
	assign w34558 = w595 ^ w597;
	assign w34709 = w34724 ^ w44827;
	assign w34675 = w34720 ^ w34709;
	assign w34672 = ~w34675;
	assign w34669 = w34725 ^ w34709;
	assign w48236 = w34698 ^ w34669;
	assign w503 = w1237 ^ w48236;
	assign w534 = w1268 ^ w503;
	assign w566 = w1300 ^ w534;
	assign w598 = w1332 ^ w566;
	assign w34644 = w595 ^ w598;
	assign w34636 = w34555 ^ w34644;
	assign w34645 = w598 ^ w592;
	assign w44828 = w34729 ^ w34731;
	assign w34687 = w44828 ^ w34684;
	assign w34784 = w34686 ^ w34687;
	assign w48229 = ~w34784;
	assign w496 = w1230 ^ w48229;
	assign w527 = w1261 ^ w496;
	assign w559 = w1293 ^ w527;
	assign w591 = w1325 ^ w559;
	assign w34562 = w591 ^ w597;
	assign w34635 = w591 ^ w34636;
	assign w34674 = w34678 ^ w44828;
	assign w34677 = w34716 ^ w34674;
	assign w34781 = w34676 ^ w34677;
	assign w34673 = w34697 ^ w34674;
	assign w48231 = w34672 ^ w34673;
	assign w48234 = ~w34781;
	assign w501 = w1235 ^ w48234;
	assign w498 = w1232 ^ w48231;
	assign w529 = w1263 ^ w498;
	assign w561 = w1295 ^ w529;
	assign w532 = w1266 ^ w501;
	assign w564 = w1298 ^ w532;
	assign w593 = w1327 ^ w561;
	assign w34557 = w593 ^ w34555;
	assign w34633 = w597 ^ w34557;
	assign w34632 = w34562 ^ w34557;
	assign w34572 = w592 ^ w593;
	assign w34640 = w34644 ^ w34572;
	assign w34646 = w593 ^ w595;
	assign w34532 = w594 ^ w593;
	assign w34643 = w598 ^ w593;
	assign w34629 = w34636 & w34640;
	assign w34561 = w34629 ^ w34558;
	assign w34623 = w34644 & w34633;
	assign w34559 = w34623 ^ w34557;
	assign w34565 = w34561 ^ w34559;
	assign w34570 = w598 ^ w34565;
	assign w596 = w1330 ^ w564;
	assign w34630 = w596 ^ w34557;
	assign w34556 = w596 ^ w598;
	assign w34631 = w34556 ^ w34646;
	assign w34639 = w34556 ^ w34562;
	assign w34637 = w34572 ^ w34639;
	assign w34642 = w596 ^ w34562;
	assign w34638 = w592 ^ w34642;
	assign w34518 = w34558 ^ w34556;
	assign w34634 = w34555 ^ w34518;
	assign w34517 = w34558 ^ w596;
	assign w34641 = w591 ^ w34517;
	assign w34628 = w34637 & w34635;
	assign w34627 = w591 & w34641;
	assign w34626 = w34645 & w34630;
	assign w34560 = w34626 ^ w34556;
	assign w34625 = w34642 & w34638;
	assign w34624 = w34639 & w34632;
	assign w34622 = w34646 & w34631;
	assign w34579 = w34622 ^ w34628;
	assign w34620 = w34579 ^ w34570;
	assign w34531 = w34622 ^ w34623;
	assign w34578 = w34531 ^ w34532;
	assign w34577 = w34578 ^ w34560;
	assign w34619 = w34625 ^ w34577;
	assign w34621 = w34643 & w34634;
	assign w34616 = w34620 & w34619;
	assign w44817 = w34621 ^ w34627;
	assign w34533 = w34565 ^ w44817;
	assign w34576 = w596 ^ w34533;
	assign w34611 = w34616 ^ w34576;
	assign w34571 = w44817 ^ w34556;
	assign w34617 = w34579 ^ w34571;
	assign w44818 = w34621 ^ w34624;
	assign w34574 = w34622 ^ w44818;
	assign w34530 = w34625 ^ w34574;
	assign w34612 = w592 ^ w34530;
	assign w34610 = w34611 & w34612;
	assign w34608 = w34616 ^ w34610;
	assign w34529 = w34610 ^ w34574;
	assign w34528 = w34610 ^ w34627;
	assign w34523 = w34528 ^ w34624;
	assign w34534 = w34560 ^ w44818;
	assign w34618 = w34534 ^ w34559;
	assign w34609 = w34610 ^ w34618;
	assign w34615 = w34616 ^ w34618;
	assign w34614 = w34617 & w34615;
	assign w34613 = w34614 ^ w34576;
	assign w34525 = w34614 ^ w34626;
	assign w34521 = w34525 ^ w34561;
	assign w34524 = w598 ^ w34521;
	assign w34601 = w34523 ^ w34524;
	assign w34522 = w34614 ^ w34570;
	assign w34520 = w596 ^ w34521;
	assign w34607 = w34618 & w34608;
	assign w34605 = w34607 ^ w34615;
	assign w34604 = w34613 & w34605;
	assign w34569 = w34604 ^ w34579;
	assign w34603 = w34569 ^ w34571;
	assign w34527 = w34604 ^ w34628;
	assign w34600 = w34569 ^ w34522;
	assign w34595 = w34609 & w591;
	assign w34594 = w34600 & w34630;
	assign w34593 = w34603 & w34642;
	assign w34592 = w34613 & w34632;
	assign w34536 = w34592 ^ w34593;
	assign w34591 = w34601 & w34633;
	assign w34586 = w34609 & w34641;
	assign w34585 = w34600 & w34645;
	assign w34552 = w34594 ^ w34585;
	assign w34584 = w34603 & w34638;
	assign w34554 = w34592 ^ w34584;
	assign w34583 = w34613 & w34639;
	assign w34582 = w34601 & w34644;
	assign w44820 = w34593 ^ w34594;
	assign w44822 = w34607 ^ w34625;
	assign w34599 = w44822 ^ w34577;
	assign w34597 = w34599 & w34636;
	assign w34588 = w34599 & w34640;
	assign w44821 = w34595 ^ w34597;
	assign w34566 = w592 ^ w44822;
	assign w34606 = w34566 ^ w34529;
	assign w34519 = w34566 ^ w34527;
	assign w34526 = w34556 ^ w34519;
	assign w34602 = w34523 ^ w34526;
	assign w34598 = w34519 ^ w34520;
	assign w34596 = w34606 & w34635;
	assign w34590 = w34598 & w34631;
	assign w34575 = w34590 ^ w44820;
	assign w34551 = w34590 ^ w34593;
	assign w34548 = ~w34551;
	assign w34547 = w34590 ^ w34591;
	assign w34541 = w34586 ^ w34575;
	assign w34538 = ~w34541;
	assign w34535 = w34591 ^ w34575;
	assign w34589 = w34602 & w34634;
	assign w34567 = w34585 ^ w34589;
	assign w34545 = ~w34567;
	assign w34544 = w34545 ^ w34583;
	assign w34540 = w34544 ^ w44821;
	assign w34543 = w34582 ^ w34540;
	assign w34587 = w34606 & w34637;
	assign w34581 = w34598 & w34646;
	assign w34580 = w34602 & w34643;
	assign w34546 = w34591 ^ w34580;
	assign w34542 = ~w34546;
	assign w34647 = w34542 ^ w34543;
	assign w48266 = ~w34647;
	assign w628 = w1362 ^ w48266;
	assign w660 = w405 ^ w628;
	assign w692 = w437 ^ w660;
	assign w724 = w469 ^ w692;
	assign w44819 = w34581 ^ w34582;
	assign w34563 = w34587 ^ w44819;
	assign w34564 = w34588 ^ w34563;
	assign w34568 = w34596 ^ w34564;
	assign w34573 = w34597 ^ w34568;
	assign w48265 = w44820 ^ w34573;
	assign w34648 = w34573 ^ w34547;
	assign w34539 = w34563 ^ w34540;
	assign w48263 = w34538 ^ w34539;
	assign w34537 = w34595 ^ w34568;
	assign w48264 = w34536 ^ w34537;
	assign w626 = w1360 ^ w48264;
	assign w658 = w403 ^ w626;
	assign w48268 = w34564 ^ w34535;
	assign w48267 = ~w34648;
	assign w627 = w1361 ^ w48265;
	assign w690 = w435 ^ w658;
	assign w722 = w467 ^ w690;
	assign w630 = w1364 ^ w48268;
	assign w662 = w407 ^ w630;
	assign w694 = w439 ^ w662;
	assign w726 = w471 ^ w694;
	assign w629 = w1363 ^ w48267;
	assign w625 = w1359 ^ w48263;
	assign w657 = w402 ^ w625;
	assign w689 = w434 ^ w657;
	assign w721 = w466 ^ w689;
	assign w661 = w406 ^ w629;
	assign w693 = w438 ^ w661;
	assign w725 = w470 ^ w693;
	assign w659 = w404 ^ w627;
	assign w691 = w436 ^ w659;
	assign w723 = w468 ^ w691;
	assign w38710 = w724 ^ w726;
	assign w38712 = w723 ^ w725;
	assign w38798 = w723 ^ w726;
	assign w38800 = w721 ^ w723;
	assign w38785 = w38710 ^ w38800;
	assign w38686 = w722 ^ w721;
	assign w38672 = w38712 ^ w38710;
	assign w38671 = w38712 ^ w724;
	assign w38797 = w726 ^ w721;
	assign w38776 = w38800 & w38785;
	assign w34550 = w34554 ^ w44819;
	assign w34553 = w44821 ^ w34550;
	assign w34650 = w34552 ^ w34553;
	assign w34549 = w34545 ^ w34550;
	assign w34649 = w34548 ^ w34549;
	assign w48261 = ~w34650;
	assign w48262 = ~w34649;
	assign w623 = w1357 ^ w48261;
	assign w655 = w400 ^ w623;
	assign w687 = w432 ^ w655;
	assign w719 = w464 ^ w687;
	assign w38716 = w719 ^ w725;
	assign w38793 = w38710 ^ w38716;
	assign w38796 = w724 ^ w38716;
	assign w38795 = w719 ^ w38671;
	assign w38781 = w719 & w38795;
	assign w43742 = w5104 ^ w5107;
	assign w5016 = w5042 ^ w43742;
	assign w5101 = w5016 ^ w5041;
	assign w5098 = w5099 ^ w5101;
	assign w5056 = w5105 ^ w43742;
	assign w5012 = w5108 ^ w5056;
	assign w5095 = w712 ^ w5012;
	assign w43741 = w5104 ^ w5110;
	assign w5053 = w43741 ^ w5038;
	assign w5100 = w5061 ^ w5053;
	assign w5097 = w5100 & w5098;
	assign w5007 = w5097 ^ w5109;
	assign w5003 = w5007 ^ w5043;
	assign w5004 = w5097 ^ w5052;
	assign w5002 = w716 ^ w5003;
	assign w5006 = w718 ^ w5003;
	assign w5015 = w5047 ^ w43741;
	assign w5058 = w716 ^ w5015;
	assign w5096 = w5097 ^ w5058;
	assign w5075 = w5096 & w5115;
	assign w5066 = w5096 & w5122;
	assign w5094 = w5099 ^ w5058;
	assign w5093 = w5094 & w5095;
	assign w5010 = w5093 ^ w5110;
	assign w5011 = w5093 ^ w5056;
	assign w5005 = w5010 ^ w5107;
	assign w5084 = w5005 ^ w5006;
	assign w5074 = w5084 & w5116;
	assign w5065 = w5084 & w5127;
	assign w5092 = w5093 ^ w5101;
	assign w5069 = w5092 & w5124;
	assign w5078 = w5092 & w711;
	assign w5091 = w5099 ^ w5093;
	assign w5090 = w5101 & w5091;
	assign w5088 = w5090 ^ w5098;
	assign w5087 = w5096 & w5088;
	assign w5051 = w5087 ^ w5061;
	assign w5083 = w5051 ^ w5004;
	assign w5009 = w5087 ^ w5111;
	assign w5077 = w5083 & w5113;
	assign w5086 = w5051 ^ w5053;
	assign w5076 = w5086 & w5125;
	assign w5067 = w5086 & w5121;
	assign w5036 = w5075 ^ w5067;
	assign w5018 = w5075 ^ w5076;
	assign w43743 = w5076 ^ w5077;
	assign w43745 = w5090 ^ w5108;
	assign w5082 = w43745 ^ w5059;
	assign w5080 = w5082 & w5119;
	assign w5071 = w5082 & w5123;
	assign w43744 = w5078 ^ w5080;
	assign w5048 = w712 ^ w43745;
	assign w5001 = w5048 ^ w5009;
	assign w5008 = w5038 ^ w5001;
	assign w5081 = w5001 ^ w5002;
	assign w5073 = w5081 & w5114;
	assign w5029 = w5073 ^ w5074;
	assign w5033 = w5073 ^ w5076;
	assign w5089 = w5048 ^ w5011;
	assign w5079 = w5089 & w5118;
	assign w5070 = w5089 & w5120;
	assign w5064 = w5081 & w5129;
	assign w5057 = w5073 ^ w43743;
	assign w5017 = w5074 ^ w5057;
	assign w5023 = w5069 ^ w5057;
	assign w5062 = w5064 ^ w5065;
	assign w5032 = w5036 ^ w5062;
	assign w5035 = w43744 ^ w5032;
	assign w5045 = w5070 ^ w5062;
	assign w5046 = w5071 ^ w5045;
	assign w5050 = w5079 ^ w5046;
	assign w5055 = w5080 ^ w5050;
	assign w48300 = w5046 ^ w5017;
	assign w5131 = w5055 ^ w5029;
	assign w48299 = ~w5131;
	assign w5019 = w5078 ^ w5050;
	assign w48296 = w5018 ^ w5019;
	assign w5030 = ~w5033;
	assign w5085 = w5005 ^ w5008;
	assign w5063 = w5085 & w5126;
	assign w5072 = w5085 & w5117;
	assign w5028 = w5074 ^ w5063;
	assign w5024 = ~w5028;
	assign w758 = w503 ^ w48300;
	assign w757 = w502 ^ w48299;
	assign w754 = w499 ^ w48296;
	assign w786 = w530 ^ w754;
	assign w789 = w533 ^ w757;
	assign w821 = w565 ^ w789;
	assign w853 = w597 ^ w821;
	assign w818 = w562 ^ w786;
	assign w850 = w594 ^ w818;
	assign w790 = w534 ^ w758;
	assign w822 = w566 ^ w790;
	assign w854 = w598 ^ w822;
	assign w48297 = w43743 ^ w5055;
	assign w755 = w500 ^ w48297;
	assign w787 = w531 ^ w755;
	assign w819 = w563 ^ w787;
	assign w851 = w595 ^ w819;
	assign w5068 = w5083 & w5128;
	assign w5034 = w5077 ^ w5068;
	assign w5133 = w5034 ^ w5035;
	assign w48293 = ~w5133;
	assign w5049 = w5068 ^ w5072;
	assign w5027 = ~w5049;
	assign w5026 = w5027 ^ w5066;
	assign w5031 = w5027 ^ w5032;
	assign w5132 = w5030 ^ w5031;
	assign w5022 = w5026 ^ w43744;
	assign w5025 = w5065 ^ w5022;
	assign w5130 = w5024 ^ w5025;
	assign w48294 = ~w5132;
	assign w48298 = ~w5130;
	assign w5021 = w5045 ^ w5022;
	assign w752 = w497 ^ w48294;
	assign w784 = w528 ^ w752;
	assign w751 = w496 ^ w48293;
	assign w783 = w527 ^ w751;
	assign w756 = w501 ^ w48298;
	assign w815 = w559 ^ w783;
	assign w847 = w591 ^ w815;
	assign w788 = w532 ^ w756;
	assign w820 = w564 ^ w788;
	assign w852 = w596 ^ w820;
	assign w816 = w560 ^ w784;
	assign w848 = w592 ^ w816;
	assign w5020 = ~w5023;
	assign w48295 = w5020 ^ w5021;
	assign w753 = w498 ^ w48295;
	assign w785 = w529 ^ w753;
	assign w817 = w561 ^ w785;
	assign w849 = w593 ^ w817;
	assign w809 = w553 ^ w777;
	assign w841 = w585 ^ w809;
	assign w624 = w1358 ^ w48262;
	assign w656 = w401 ^ w624;
	assign w688 = w433 ^ w656;
	assign w720 = w465 ^ w688;
	assign w38709 = w720 ^ w722;
	assign w38711 = w721 ^ w38709;
	assign w38787 = w725 ^ w38711;
	assign w38784 = w724 ^ w38711;
	assign w38786 = w38716 ^ w38711;
	assign w38792 = w720 ^ w38796;
	assign w38790 = w38709 ^ w38798;
	assign w38789 = w719 ^ w38790;
	assign w38726 = w720 ^ w721;
	assign w38791 = w38726 ^ w38793;
	assign w38794 = w38798 ^ w38726;
	assign w38788 = w38709 ^ w38672;
	assign w38799 = w726 ^ w720;
	assign w38783 = w38790 & w38794;
	assign w38715 = w38783 ^ w38712;
	assign w38782 = w38791 & w38789;
	assign w38733 = w38776 ^ w38782;
	assign w38780 = w38799 & w38784;
	assign w38714 = w38780 ^ w38710;
	assign w38779 = w38796 & w38792;
	assign w38778 = w38793 & w38786;
	assign w38777 = w38798 & w38787;
	assign w38713 = w38777 ^ w38711;
	assign w38719 = w38715 ^ w38713;
	assign w38724 = w726 ^ w38719;
	assign w38774 = w38733 ^ w38724;
	assign w38685 = w38776 ^ w38777;
	assign w38732 = w38685 ^ w38686;
	assign w38731 = w38732 ^ w38714;
	assign w38773 = w38779 ^ w38731;
	assign w38775 = w38797 & w38788;
	assign w38770 = w38774 & w38773;
	assign w812 = w556 ^ w780;
	assign w844 = w588 ^ w812;
	assign w44993 = w38775 ^ w38781;
	assign w38725 = w44993 ^ w38710;
	assign w38771 = w38733 ^ w38725;
	assign w38687 = w38719 ^ w44993;
	assign w38730 = w724 ^ w38687;
	assign w38765 = w38770 ^ w38730;
	assign w44994 = w38775 ^ w38778;
	assign w38728 = w38776 ^ w44994;
	assign w38684 = w38779 ^ w38728;
	assign w38766 = w720 ^ w38684;
	assign w38764 = w38765 & w38766;
	assign w38762 = w38770 ^ w38764;
	assign w38683 = w38764 ^ w38728;
	assign w38682 = w38764 ^ w38781;
	assign w38677 = w38682 ^ w38778;
	assign w38688 = w38714 ^ w44994;
	assign w38772 = w38688 ^ w38713;
	assign w38763 = w38764 ^ w38772;
	assign w38769 = w38770 ^ w38772;
	assign w38768 = w38771 & w38769;
	assign w38767 = w38768 ^ w38730;
	assign w38679 = w38768 ^ w38780;
	assign w38675 = w38679 ^ w38715;
	assign w38678 = w726 ^ w38675;
	assign w38755 = w38677 ^ w38678;
	assign w38676 = w38768 ^ w38724;
	assign w38674 = w724 ^ w38675;
	assign w38761 = w38772 & w38762;
	assign w38759 = w38761 ^ w38769;
	assign w38758 = w38767 & w38759;
	assign w38723 = w38758 ^ w38733;
	assign w38757 = w38723 ^ w38725;
	assign w38681 = w38758 ^ w38782;
	assign w38754 = w38723 ^ w38676;
	assign w38749 = w38763 & w719;
	assign w38748 = w38754 & w38784;
	assign w38747 = w38757 & w38796;
	assign w38746 = w38767 & w38786;
	assign w38690 = w38746 ^ w38747;
	assign w38745 = w38755 & w38787;
	assign w38740 = w38763 & w38795;
	assign w38739 = w38754 & w38799;
	assign w38706 = w38748 ^ w38739;
	assign w38738 = w38757 & w38792;
	assign w38708 = w38746 ^ w38738;
	assign w38737 = w38767 & w38793;
	assign w38736 = w38755 & w38798;
	assign w44995 = w38747 ^ w38748;
	assign w44997 = w38761 ^ w38779;
	assign w38720 = w720 ^ w44997;
	assign w38760 = w38720 ^ w38683;
	assign w38750 = w38760 & w38789;
	assign w38741 = w38760 & w38791;
	assign w38673 = w38720 ^ w38681;
	assign w38752 = w38673 ^ w38674;
	assign w38744 = w38752 & w38785;
	assign w38705 = w38744 ^ w38747;
	assign w38702 = ~w38705;
	assign w38701 = w38744 ^ w38745;
	assign w38735 = w38752 & w38800;
	assign w43606 = w38735 ^ w38736;
	assign w38704 = w38708 ^ w43606;
	assign w38717 = w38741 ^ w43606;
	assign w38680 = w38710 ^ w38673;
	assign w38729 = w38744 ^ w44995;
	assign w38695 = w38740 ^ w38729;
	assign w38692 = ~w38695;
	assign w38689 = w38745 ^ w38729;
	assign w38756 = w38677 ^ w38680;
	assign w38734 = w38756 & w38797;
	assign w38700 = w38745 ^ w38734;
	assign w38696 = ~w38700;
	assign w38743 = w38756 & w38788;
	assign w38721 = w38739 ^ w38743;
	assign w38699 = ~w38721;
	assign w38703 = w38699 ^ w38704;
	assign w38803 = w38702 ^ w38703;
	assign w48302 = ~w38803;
	assign w760 = w505 ^ w48302;
	assign w792 = w536 ^ w760;
	assign w824 = w568 ^ w792;
	assign w856 = w600 ^ w824;
	assign w38698 = w38699 ^ w38737;
	assign w38753 = w44997 ^ w38731;
	assign w38751 = w38753 & w38790;
	assign w38742 = w38753 & w38794;
	assign w38718 = w38742 ^ w38717;
	assign w38722 = w38750 ^ w38718;
	assign w38727 = w38751 ^ w38722;
	assign w48305 = w44995 ^ w38727;
	assign w763 = w508 ^ w48305;
	assign w795 = w539 ^ w763;
	assign w38802 = w38727 ^ w38701;
	assign w38691 = w38749 ^ w38722;
	assign w48304 = w38690 ^ w38691;
	assign w762 = w507 ^ w48304;
	assign w794 = w538 ^ w762;
	assign w826 = w570 ^ w794;
	assign w858 = w602 ^ w826;
	assign w48308 = w38718 ^ w38689;
	assign w48307 = ~w38802;
	assign w827 = w571 ^ w795;
	assign w766 = w510 ^ w48308;
	assign w798 = w542 ^ w766;
	assign w2048 = w509 ^ w48307;
	assign w765 = ~w2048;
	assign w797 = w541 ^ w765;
	assign w829 = w573 ^ w797;
	assign w861 = w605 ^ w829;
	assign w830 = w574 ^ w798;
	assign w862 = w606 ^ w830;
	assign w859 = w603 ^ w827;
	assign w44996 = w38749 ^ w38751;
	assign w38707 = w44996 ^ w38704;
	assign w38804 = w38706 ^ w38707;
	assign w48301 = ~w38804;
	assign w759 = w504 ^ w48301;
	assign w791 = w535 ^ w759;
	assign w823 = w567 ^ w791;
	assign w855 = w599 ^ w823;
	assign w38694 = w38698 ^ w44996;
	assign w38697 = w38736 ^ w38694;
	assign w38801 = w38696 ^ w38697;
	assign w38693 = w38717 ^ w38694;
	assign w48303 = w38692 ^ w38693;
	assign w761 = w506 ^ w48303;
	assign w793 = w537 ^ w761;
	assign w825 = w569 ^ w793;
	assign w857 = w601 ^ w825;
	assign w48306 = ~w38801;
	assign w764 = w45168 ^ w48306;
	assign w796 = w540 ^ w764;
	assign w828 = w572 ^ w796;
	assign w860 = w604 ^ w828;
	assign w44998 = w38909 ^ w38915;
	assign w38821 = w38853 ^ w44998;
	assign w38864 = w604 ^ w38821;
	assign w38899 = w38904 ^ w38864;
	assign w38859 = w44998 ^ w38844;
	assign w38905 = w38867 ^ w38859;
	assign w44999 = w38909 ^ w38912;
	assign w38862 = w38910 ^ w44999;
	assign w38818 = w38913 ^ w38862;
	assign w38900 = w600 ^ w38818;
	assign w38898 = w38899 & w38900;
	assign w38817 = w38898 ^ w38862;
	assign w38896 = w38904 ^ w38898;
	assign w38816 = w38898 ^ w38915;
	assign w38811 = w38816 ^ w38912;
	assign w38822 = w38848 ^ w44999;
	assign w38906 = w38822 ^ w38847;
	assign w38897 = w38898 ^ w38906;
	assign w38903 = w38904 ^ w38906;
	assign w38902 = w38905 & w38903;
	assign w38901 = w38902 ^ w38864;
	assign w38813 = w38902 ^ w38914;
	assign w38809 = w38813 ^ w38849;
	assign w38812 = w606 ^ w38809;
	assign w38889 = w38811 ^ w38812;
	assign w38810 = w38902 ^ w38858;
	assign w38808 = w604 ^ w38809;
	assign w38895 = w38906 & w38896;
	assign w38893 = w38895 ^ w38903;
	assign w38892 = w38901 & w38893;
	assign w38857 = w38892 ^ w38867;
	assign w38891 = w38857 ^ w38859;
	assign w38815 = w38892 ^ w38916;
	assign w38888 = w38857 ^ w38810;
	assign w38883 = w38897 & w599;
	assign w38882 = w38888 & w38918;
	assign w38881 = w38891 & w38930;
	assign w38880 = w38901 & w38920;
	assign w38824 = w38880 ^ w38881;
	assign w38879 = w38889 & w38921;
	assign w38874 = w38897 & w38929;
	assign w38873 = w38888 & w38933;
	assign w38840 = w38882 ^ w38873;
	assign w38872 = w38891 & w38926;
	assign w38842 = w38880 ^ w38872;
	assign w38871 = w38901 & w38927;
	assign w38870 = w38889 & w38932;
	assign w45001 = w38881 ^ w38882;
	assign w45003 = w38895 ^ w38913;
	assign w38887 = w45003 ^ w38865;
	assign w38885 = w38887 & w38924;
	assign w45002 = w38883 ^ w38885;
	assign w38876 = w38887 & w38928;
	assign w38854 = w600 ^ w45003;
	assign w38894 = w38854 ^ w38817;
	assign w38807 = w38854 ^ w38815;
	assign w38814 = w38844 ^ w38807;
	assign w38890 = w38811 ^ w38814;
	assign w38886 = w38807 ^ w38808;
	assign w38884 = w38894 & w38923;
	assign w38878 = w38886 & w38919;
	assign w38863 = w38878 ^ w45001;
	assign w38839 = w38878 ^ w38881;
	assign w38836 = ~w38839;
	assign w38835 = w38878 ^ w38879;
	assign w38829 = w38874 ^ w38863;
	assign w38826 = ~w38829;
	assign w38823 = w38879 ^ w38863;
	assign w38877 = w38890 & w38922;
	assign w38855 = w38873 ^ w38877;
	assign w38833 = ~w38855;
	assign w38832 = w38833 ^ w38871;
	assign w38828 = w38832 ^ w45002;
	assign w38831 = w38870 ^ w38828;
	assign w38875 = w38894 & w38925;
	assign w38869 = w38886 & w38934;
	assign w38868 = w38890 & w38931;
	assign w38834 = w38879 ^ w38868;
	assign w38830 = ~w38834;
	assign w38935 = w38830 ^ w38831;
	assign w48274 = ~w38935;
	assign w636 = w1370 ^ w48274;
	assign w668 = w413 ^ w636;
	assign w700 = w445 ^ w668;
	assign w732 = w477 ^ w700;
	assign w45000 = w38869 ^ w38870;
	assign w38851 = w38875 ^ w45000;
	assign w38852 = w38876 ^ w38851;
	assign w48276 = w38852 ^ w38823;
	assign w38856 = w38884 ^ w38852;
	assign w38825 = w38883 ^ w38856;
	assign w48272 = w38824 ^ w38825;
	assign w634 = w1368 ^ w48272;
	assign w666 = w411 ^ w634;
	assign w38861 = w38885 ^ w38856;
	assign w48273 = w45001 ^ w38861;
	assign w635 = w1369 ^ w48273;
	assign w38936 = w38861 ^ w38835;
	assign w48275 = ~w38936;
	assign w637 = w1371 ^ w48275;
	assign w669 = w414 ^ w637;
	assign w701 = w446 ^ w669;
	assign w733 = w478 ^ w701;
	assign w38827 = w38851 ^ w38828;
	assign w48271 = w38826 ^ w38827;
	assign w698 = w443 ^ w666;
	assign w730 = w475 ^ w698;
	assign w638 = w1372 ^ w48276;
	assign w670 = w415 ^ w638;
	assign w702 = w447 ^ w670;
	assign w734 = w479 ^ w702;
	assign w36164 = w732 ^ w734;
	assign w667 = w412 ^ w635;
	assign w699 = w444 ^ w667;
	assign w731 = w476 ^ w699;
	assign w36166 = w731 ^ w733;
	assign w36252 = w731 ^ w734;
	assign w36126 = w36166 ^ w36164;
	assign w36125 = w36166 ^ w732;
	assign w633 = w1367 ^ w48271;
	assign w665 = w410 ^ w633;
	assign w697 = w442 ^ w665;
	assign w729 = w474 ^ w697;
	assign w36254 = w729 ^ w731;
	assign w36239 = w36164 ^ w36254;
	assign w36251 = w734 ^ w729;
	assign w36230 = w36254 & w36239;
	assign w36140 = w730 ^ w729;
	assign w38838 = w38842 ^ w45000;
	assign w38841 = w45002 ^ w38838;
	assign w38938 = w38840 ^ w38841;
	assign w38837 = w38833 ^ w38838;
	assign w38937 = w38836 ^ w38837;
	assign w48269 = ~w38938;
	assign w631 = w1365 ^ w48269;
	assign w663 = w408 ^ w631;
	assign w48270 = ~w38937;
	assign w632 = w1366 ^ w48270;
	assign w664 = w409 ^ w632;
	assign w696 = w441 ^ w664;
	assign w728 = w473 ^ w696;
	assign w36163 = w728 ^ w730;
	assign w36165 = w729 ^ w36163;
	assign w36241 = w733 ^ w36165;
	assign w36238 = w732 ^ w36165;
	assign w36244 = w36163 ^ w36252;
	assign w36180 = w728 ^ w729;
	assign w36248 = w36252 ^ w36180;
	assign w36242 = w36163 ^ w36126;
	assign w36253 = w734 ^ w728;
	assign w36237 = w36244 & w36248;
	assign w36169 = w36237 ^ w36166;
	assign w36234 = w36253 & w36238;
	assign w36168 = w36234 ^ w36164;
	assign w36231 = w36252 & w36241;
	assign w36167 = w36231 ^ w36165;
	assign w36173 = w36169 ^ w36167;
	assign w36178 = w734 ^ w36173;
	assign w36139 = w36230 ^ w36231;
	assign w36186 = w36139 ^ w36140;
	assign w36185 = w36186 ^ w36168;
	assign w36229 = w36251 & w36242;
	assign w695 = w440 ^ w663;
	assign w727 = w472 ^ w695;
	assign w36243 = w727 ^ w36244;
	assign w36170 = w727 ^ w733;
	assign w36240 = w36170 ^ w36165;
	assign w36247 = w36164 ^ w36170;
	assign w36245 = w36180 ^ w36247;
	assign w36250 = w732 ^ w36170;
	assign w36246 = w728 ^ w36250;
	assign w36249 = w727 ^ w36125;
	assign w36236 = w36245 & w36243;
	assign w36187 = w36230 ^ w36236;
	assign w36228 = w36187 ^ w36178;
	assign w36235 = w36249 & w727;
	assign w36233 = w36250 & w36246;
	assign w36227 = w36233 ^ w36185;
	assign w36232 = w36247 & w36240;
	assign w36224 = w36228 & w36227;
	assign w44885 = w36229 ^ w36235;
	assign w36141 = w36173 ^ w44885;
	assign w36184 = w732 ^ w36141;
	assign w36219 = w36224 ^ w36184;
	assign w36179 = w44885 ^ w36164;
	assign w36225 = w36187 ^ w36179;
	assign w44886 = w36229 ^ w36232;
	assign w36182 = w36230 ^ w44886;
	assign w36138 = w36233 ^ w36182;
	assign w36220 = w728 ^ w36138;
	assign w36218 = w36219 & w36220;
	assign w36216 = w36224 ^ w36218;
	assign w36137 = w36218 ^ w36182;
	assign w36136 = w36218 ^ w36235;
	assign w36131 = w36136 ^ w36232;
	assign w36142 = w36168 ^ w44886;
	assign w36226 = w36142 ^ w36167;
	assign w36217 = w36218 ^ w36226;
	assign w36223 = w36224 ^ w36226;
	assign w36222 = w36225 & w36223;
	assign w36221 = w36222 ^ w36184;
	assign w36133 = w36222 ^ w36234;
	assign w36129 = w36133 ^ w36169;
	assign w36132 = w734 ^ w36129;
	assign w36209 = w36131 ^ w36132;
	assign w36130 = w36222 ^ w36178;
	assign w36128 = w732 ^ w36129;
	assign w36215 = w36226 & w36216;
	assign w36213 = w36215 ^ w36223;
	assign w36212 = w36221 & w36213;
	assign w36177 = w36212 ^ w36187;
	assign w36211 = w36177 ^ w36179;
	assign w36135 = w36212 ^ w36236;
	assign w36208 = w36177 ^ w36130;
	assign w36203 = w36217 & w727;
	assign w36202 = w36208 & w36238;
	assign w36201 = w36211 & w36250;
	assign w36200 = w36221 & w36240;
	assign w36144 = w36200 ^ w36201;
	assign w36199 = w36209 & w36241;
	assign w36194 = w36217 & w36249;
	assign w36193 = w36208 & w36253;
	assign w36160 = w36202 ^ w36193;
	assign w36192 = w36211 & w36246;
	assign w36162 = w36200 ^ w36192;
	assign w36191 = w36221 & w36247;
	assign w36190 = w36209 & w36252;
	assign w44888 = w36201 ^ w36202;
	assign w44890 = w36215 ^ w36233;
	assign w36207 = w44890 ^ w36185;
	assign w36205 = w36207 & w36244;
	assign w44889 = w36203 ^ w36205;
	assign w36196 = w36207 & w36248;
	assign w36174 = w728 ^ w44890;
	assign w36214 = w36174 ^ w36137;
	assign w36127 = w36174 ^ w36135;
	assign w36134 = w36164 ^ w36127;
	assign w36210 = w36131 ^ w36134;
	assign w36206 = w36127 ^ w36128;
	assign w36204 = w36214 & w36243;
	assign w36198 = w36206 & w36239;
	assign w36183 = w36198 ^ w44888;
	assign w36159 = w36198 ^ w36201;
	assign w36156 = ~w36159;
	assign w36155 = w36198 ^ w36199;
	assign w36149 = w36194 ^ w36183;
	assign w36146 = ~w36149;
	assign w36143 = w36199 ^ w36183;
	assign w36197 = w36210 & w36242;
	assign w36175 = w36193 ^ w36197;
	assign w36153 = ~w36175;
	assign w36152 = w36153 ^ w36191;
	assign w36148 = w36152 ^ w44889;
	assign w36151 = w36190 ^ w36148;
	assign w36195 = w36214 & w36245;
	assign w36189 = w36206 & w36254;
	assign w36188 = w36210 & w36251;
	assign w36154 = w36199 ^ w36188;
	assign w36150 = ~w36154;
	assign w36255 = w36150 ^ w36151;
	assign w48282 = ~w36255;
	assign w740 = w485 ^ w48282;
	assign w772 = w516 ^ w740;
	assign w804 = w548 ^ w772;
	assign w836 = w580 ^ w804;
	assign w44887 = w36189 ^ w36190;
	assign w36158 = w36162 ^ w44887;
	assign w36161 = w44889 ^ w36158;
	assign w36258 = w36160 ^ w36161;
	assign w36157 = w36153 ^ w36158;
	assign w36257 = w36156 ^ w36157;
	assign w48278 = ~w36257;
	assign w736 = w481 ^ w48278;
	assign w768 = w512 ^ w736;
	assign w800 = w544 ^ w768;
	assign w832 = w576 ^ w800;
	assign w48277 = ~w36258;
	assign w735 = w480 ^ w48277;
	assign w767 = w511 ^ w735;
	assign w799 = w543 ^ w767;
	assign w831 = w575 ^ w799;
	assign w36171 = w36195 ^ w44887;
	assign w36172 = w36196 ^ w36171;
	assign w36176 = w36204 ^ w36172;
	assign w36181 = w36205 ^ w36176;
	assign w48281 = w44888 ^ w36181;
	assign w36256 = w36181 ^ w36155;
	assign w36147 = w36171 ^ w36148;
	assign w48279 = w36146 ^ w36147;
	assign w36145 = w36203 ^ w36176;
	assign w48280 = w36144 ^ w36145;
	assign w48284 = w36172 ^ w36143;
	assign w48283 = ~w36256;
	assign w742 = w487 ^ w48284;
	assign w774 = w518 ^ w742;
	assign w739 = w484 ^ w48281;
	assign w771 = w515 ^ w739;
	assign w803 = w547 ^ w771;
	assign w835 = w579 ^ w803;
	assign w738 = w483 ^ w48280;
	assign w770 = w514 ^ w738;
	assign w802 = w546 ^ w770;
	assign w834 = w578 ^ w802;
	assign w806 = w550 ^ w774;
	assign w838 = w582 ^ w806;
	assign w737 = w482 ^ w48279;
	assign w769 = w513 ^ w737;
	assign w801 = w545 ^ w769;
	assign w833 = w577 ^ w801;
	assign w741 = w486 ^ w48283;
	assign w773 = w517 ^ w741;
	assign w805 = w549 ^ w773;
	assign w837 = w581 ^ w805;
	assign w776 = w520 ^ w744;
	assign w808 = w552 ^ w776;
	assign w840 = w584 ^ w808;
	assign w45172 = ~w5399;
	assign w6166 = w48469 ^ w45172;
	assign w45173 = ~w5400;
	assign w6152 = w6031 ^ w45173;
	assign w6143 = w45173 ^ w5936;
	assign w48359 = w6144 ^ w6143;
	assign w47714 = w48359 ^ w50;
	assign w21246 = w47714 ^ w47712;
	assign w21132 = w47713 ^ w47714;
	assign w45174 = ~w5401;
	assign w45175 = ~w5267;
	assign w45176 = ~w5532;
	assign w6175 = w45176 ^ w36122;
	assign w45177 = ~w5534;
	assign w6095 = w6124 ^ w45177;
	assign w6106 = w45177 ^ w29021;
	assign w48335 = w6107 ^ w6106;
	assign w47738 = w48335 ^ w26;
	assign w45178 = ~w5535;
	assign w6235 = w6028 ^ w45178;
	assign w45179 = ~w5398;
	assign w45180 = ~w5666;
	assign w6064 = w45180 ^ w48500;
	assign w45181 = ~w5667;
	assign w5969 = w48496 ^ w45181;
	assign w6058 = w5969 ^ w6034;
	assign w48420 = w48497 ^ w6058;
	assign w47653 = w48420 ^ w111;
	assign w45182 = ~w5668;
	assign w45183 = ~w5669;
	assign w45184 = ~w5800;
	assign w45185 = ~w5801;
	assign w6182 = w6032 ^ w45185;
	assign w45186 = ~w5802;
	assign w6249 = w6025 ^ w45186;
	assign w6171 = w6169 ^ w45186;
	assign w45187 = ~w5803;
	assign w6257 = w6255 ^ w45187;
	assign w45188 = ~w5934;
	assign w6118 = w45188 ^ w48459;
	assign w45189 = ~w5935;
	assign w6013 = w45189 ^ w45172;
	assign w6148 = w45189 ^ w45188;
	assign w6150 = w6013 ^ w6030;
	assign w48364 = w48473 ^ w6150;
	assign w47709 = w48364 ^ w55;
	assign w21244 = w47712 ^ w47709;
	assign w21243 = w47709 ^ w47714;
	assign w6140 = w6031 ^ w45189;
	assign w45190 = ~w5937;
	assign w6263 = w45174 ^ w45190;
	assign w45482 = ~w21517;
	assign w6282 = w6019 ^ w45482;
	assign w6224 = w45482 ^ w48498;
	assign w45483 = ~w21518;
	assign w6267 = w45483 ^ w45182;
	assign w45486 = ~w21651;
	assign w5967 = w45486 ^ w48478;
	assign w6187 = w5967 ^ w5982;
	assign w48383 = w48474 ^ w6187;
	assign w6170 = w6245 ^ w45486;
	assign w47690 = w48383 ^ w74;
	assign w48375 = w6171 ^ w6170;
	assign w47698 = w48375 ^ w66;
	assign w21112 = w47698 ^ w47696;
	assign w20998 = w47697 ^ w47698;
	assign w45487 = ~w21652;
	assign w5966 = w45487 ^ w45175;
	assign w6256 = w5266 ^ w45487;
	assign w6197 = w5966 ^ w6025;
	assign w48389 = w45187 ^ w6197;
	assign w47684 = w48389 ^ w80;
	assign w6208 = w5966 ^ w6032;
	assign w5950 = w6257 ^ w6256;
	assign w45488 = ~w21515;
	assign w6079 = w5969 ^ w45488;
	assign w45489 = ~w21516;
	assign w45490 = ~w21785;
	assign w6060 = w45490 ^ w45182;
	assign w48423 = w6061 ^ w6060;
	assign w6004 = w45490 ^ w45482;
	assign w6073 = w5994 ^ w6004;
	assign w48431 = w48502 ^ w6073;
	assign w47650 = w48423 ^ w114;
	assign w20844 = w47650 ^ w47648;
	assign w20730 = w47649 ^ w47650;
	assign w47642 = w48431 ^ w122;
	assign w32100 = w47642 ^ w47640;
	assign w45491 = ~w21786;
	assign w5984 = w45491 ^ w45483;
	assign w6223 = w5984 ^ w6022;
	assign w48405 = w45183 ^ w6223;
	assign w47668 = w48405 ^ w96;
	assign w6281 = w45491 ^ w45183;
	assign w5939 = w6282 ^ w6281;
	assign w6044 = w5984 ^ w6033;
	assign w45492 = ~w21649;
	assign w6178 = w5265 ^ w45492;
	assign w5996 = w45492 ^ w48482;
	assign w6202 = w5996 ^ w45184;
	assign w48394 = w6202 ^ w6201;
	assign w6220 = w5996 ^ w6001;
	assign w47679 = w48394 ^ w85;
	assign w45493 = ~w21650;
	assign w6003 = w45493 ^ w48483;
	assign w6194 = w6003 ^ w6032;
	assign w48388 = w48477 ^ w6194;
	assign w6181 = w48484 ^ w45493;
	assign w48380 = w6182 ^ w6181;
	assign w6203 = w6003 ^ w45185;
	assign w6205 = ~w6203;
	assign w47693 = w48380 ^ w71;
	assign w21110 = w47696 ^ w47693;
	assign w21109 = w47693 ^ w47698;
	assign w47685 = w48388 ^ w79;
	assign w6409 = w47685 ^ w47690;
	assign w45494 = ~w21919;
	assign w5978 = w45494 ^ w45186;
	assign w48374 = w5950 ^ w5978;
	assign w6185 = w5966 ^ w5978;
	assign w6213 = w5974 ^ w5978;
	assign w48399 = w48485 ^ w6213;
	assign w6199 = w45494 ^ w5266;
	assign w48391 = w6200 ^ w6199;
	assign w47682 = w48391 ^ w82;
	assign w25668 = w47682 ^ w47680;
	assign w25554 = w47681 ^ w47682;
	assign w47699 = w48374 ^ w65;
	assign w21021 = w47699 ^ w47697;
	assign w21023 = w47698 ^ w21021;
	assign w21102 = w21021 ^ w21110;
	assign w21038 = w47699 ^ w47698;
	assign w21106 = w21110 ^ w21038;
	assign w21111 = w47693 ^ w47699;
	assign w21095 = w21102 & w21106;
	assign w47674 = w48399 ^ w90;
	assign w45495 = ~w21920;
	assign w5970 = w45495 ^ w45187;
	assign w6168 = w5970 ^ w6024;
	assign w48373 = w45175 ^ w6168;
	assign w6183 = w5970 ^ w6029;
	assign w6248 = w45495 ^ w45175;
	assign w5953 = w6249 ^ w6248;
	assign w48390 = w5953 ^ w5967;
	assign w48397 = w45495 ^ w6208;
	assign w6209 = w5967 ^ w5970;
	assign w47676 = w48397 ^ w88;
	assign w47683 = w48390 ^ w81;
	assign w25577 = w47683 ^ w47681;
	assign w25579 = w47682 ^ w25577;
	assign w25652 = w47679 ^ w25579;
	assign w25594 = w47683 ^ w47682;
	assign w47700 = w48373 ^ w64;
	assign w21101 = w47700 ^ w21102;
	assign w48381 = w45487 ^ w6183;
	assign w47692 = w48381 ^ w72;
	assign w6211 = ~w6209;
	assign w45496 = ~w21783;
	assign w6009 = w45180 ^ w45496;
	assign w6077 = w6009 ^ w6017;
	assign w6066 = w5969 ^ w6009;
	assign w48427 = w45489 ^ w6066;
	assign w47646 = w48427 ^ w118;
	assign w20756 = w47648 ^ w47646;
	assign w6038 = ~w6009;
	assign w6040 = w6038 ^ w45488;
	assign w48410 = w6040 ^ w6039;
	assign w47663 = w48410 ^ w101;
	assign w45497 = ~w21784;
	assign w6078 = w45497 ^ w45496;
	assign w48435 = w6079 ^ w6078;
	assign w6067 = w45497 ^ w45181;
	assign w48428 = w6068 ^ w6067;
	assign w6011 = w45497 ^ w45489;
	assign w6080 = w6011 ^ w6033;
	assign w48436 = w48505 ^ w6080;
	assign w6056 = w6011 ^ w45180;
	assign w47645 = w48428 ^ w119;
	assign w20842 = w47648 ^ w47645;
	assign w20841 = w47645 ^ w47650;
	assign w47637 = w48436 ^ w127;
	assign w32098 = w47640 ^ w47637;
	assign w32097 = w47637 ^ w47642;
	assign w47638 = w48435 ^ w126;
	assign w32012 = w47640 ^ w47638;
	assign w45498 = ~w22053;
	assign w6053 = w45498 ^ w6231;
	assign w5965 = w45498 ^ w45177;
	assign w6112 = w5965 ^ w5988;
	assign w48311 = w48452 ^ w6112;
	assign w47762 = w48311 ^ w2;
	assign w32502 = w47762 ^ w47760;
	assign w32388 = w47761 ^ w47762;
	assign w45499 = ~w22054;
	assign w5964 = w45499 ^ w45178;
	assign w6087 = w5964 ^ w6026;
	assign w6238 = w29021 ^ w45499;
	assign w6212 = w5964 ^ w6027;
	assign w45500 = ~w21917;
	assign w6007 = w45500 ^ w45184;
	assign w6192 = w5989 ^ w6007;
	assign w6204 = w45500 ^ w5264;
	assign w48402 = w45500 ^ w6220;
	assign w48386 = w45492 ^ w6192;
	assign w48395 = w6205 ^ w6204;
	assign w6221 = w6003 ^ w6007;
	assign w47671 = w48402 ^ w93;
	assign w47678 = w48395 ^ w86;
	assign w25655 = w47678 ^ w25579;
	assign w25580 = w47680 ^ w47678;
	assign w25584 = w47684 ^ w47678;
	assign w25654 = w25584 ^ w25579;
	assign w25664 = w47679 ^ w25584;
	assign w25660 = w47683 ^ w25664;
	assign w25539 = w25580 ^ w47679;
	assign w25663 = w47684 ^ w25539;
	assign w25649 = w47684 & w25663;
	assign w25647 = w25664 & w25660;
	assign w47687 = w48386 ^ w77;
	assign w6322 = w47687 ^ w47685;
	assign w6172 = w6007 ^ w48491;
	assign w6174 = ~w6172;
	assign w48378 = w6174 ^ w6173;
	assign w47695 = w48378 ^ w69;
	assign w21096 = w47695 ^ w21023;
	assign w21022 = w47695 ^ w47693;
	assign w21097 = w21022 ^ w21112;
	assign w21092 = w21111 & w21096;
	assign w21026 = w21092 ^ w21022;
	assign w21088 = w21112 & w21097;
	assign w45501 = ~w21918;
	assign w6018 = w45501 ^ w45185;
	assign w48403 = w45501 ^ w6221;
	assign w6222 = w6018 ^ w6029;
	assign w48404 = w48488 ^ w6222;
	assign w6179 = w6018 ^ w45184;
	assign w6180 = w6179 ^ w6178;
	assign w48379 = ~w6180;
	assign w6193 = w5996 ^ w6018;
	assign w48387 = w45493 ^ w6193;
	assign w6206 = w45501 ^ w5265;
	assign w47694 = w48379 ^ w70;
	assign w21099 = w47694 ^ w21023;
	assign w21024 = w47696 ^ w47694;
	assign w21027 = w21095 ^ w21024;
	assign w21028 = w47700 ^ w47694;
	assign w21098 = w21028 ^ w21023;
	assign w21105 = w21022 ^ w21028;
	assign w21103 = w21038 ^ w21105;
	assign w21108 = w47695 ^ w21028;
	assign w21104 = w47699 ^ w21108;
	assign w20984 = w21024 ^ w21022;
	assign w21100 = w21021 ^ w20984;
	assign w20983 = w21024 ^ w47695;
	assign w21107 = w47700 ^ w20983;
	assign w21094 = w21103 & w21101;
	assign w21045 = w21088 ^ w21094;
	assign w21093 = w47700 & w21107;
	assign w21091 = w21108 & w21104;
	assign w21090 = w21105 & w21098;
	assign w21089 = w21110 & w21099;
	assign w21025 = w21089 ^ w21023;
	assign w21031 = w21027 ^ w21025;
	assign w21036 = w47693 ^ w21031;
	assign w21086 = w21045 ^ w21036;
	assign w20997 = w21088 ^ w21089;
	assign w21044 = w20997 ^ w20998;
	assign w21043 = w21044 ^ w21026;
	assign w21085 = w21091 ^ w21043;
	assign w21087 = w21109 & w21100;
	assign w21082 = w21086 & w21085;
	assign w47686 = w48387 ^ w78;
	assign w6328 = w47692 ^ w47686;
	assign w6408 = w47687 ^ w6328;
	assign w6405 = w6322 ^ w6328;
	assign w47670 = w48403 ^ w94;
	assign w32150 = w47676 ^ w47670;
	assign w32230 = w47671 ^ w32150;
	assign w47669 = w48404 ^ w95;
	assign w32144 = w47671 ^ w47669;
	assign w32227 = w32144 ^ w32150;
	assign w32231 = w47669 ^ w47674;
	assign w44249 = w21087 ^ w21093;
	assign w20999 = w21031 ^ w44249;
	assign w21042 = w47695 ^ w20999;
	assign w21077 = w21082 ^ w21042;
	assign w21037 = w44249 ^ w21022;
	assign w21083 = w21045 ^ w21037;
	assign w44250 = w21087 ^ w21090;
	assign w21040 = w21088 ^ w44250;
	assign w20996 = w21091 ^ w21040;
	assign w21078 = w47699 ^ w20996;
	assign w21076 = w21077 & w21078;
	assign w20995 = w21076 ^ w21040;
	assign w21074 = w21082 ^ w21076;
	assign w20994 = w21076 ^ w21093;
	assign w20989 = w20994 ^ w21090;
	assign w21000 = w21026 ^ w44250;
	assign w21084 = w21000 ^ w21025;
	assign w21075 = w21076 ^ w21084;
	assign w21081 = w21082 ^ w21084;
	assign w21080 = w21083 & w21081;
	assign w21079 = w21080 ^ w21042;
	assign w20991 = w21080 ^ w21092;
	assign w20987 = w20991 ^ w21027;
	assign w20990 = w47693 ^ w20987;
	assign w21067 = w20989 ^ w20990;
	assign w20988 = w21080 ^ w21036;
	assign w20986 = w47695 ^ w20987;
	assign w21073 = w21084 & w21074;
	assign w21071 = w21073 ^ w21081;
	assign w21070 = w21079 & w21071;
	assign w21035 = w21070 ^ w21045;
	assign w21069 = w21035 ^ w21037;
	assign w20993 = w21070 ^ w21094;
	assign w21066 = w21035 ^ w20988;
	assign w21061 = w21075 & w47700;
	assign w21060 = w21066 & w21096;
	assign w21059 = w21069 & w21108;
	assign w21058 = w21079 & w21098;
	assign w21002 = w21058 ^ w21059;
	assign w21057 = w21067 & w21099;
	assign w21052 = w21075 & w21107;
	assign w21051 = w21066 & w21111;
	assign w21018 = w21060 ^ w21051;
	assign w21050 = w21069 & w21104;
	assign w21020 = w21058 ^ w21050;
	assign w21049 = w21079 & w21105;
	assign w21048 = w21067 & w21110;
	assign w44252 = w21059 ^ w21060;
	assign w44254 = w21073 ^ w21091;
	assign w21065 = w44254 ^ w21043;
	assign w21063 = w21065 & w21102;
	assign w44253 = w21061 ^ w21063;
	assign w21054 = w21065 & w21106;
	assign w21032 = w47699 ^ w44254;
	assign w21072 = w21032 ^ w20995;
	assign w20985 = w21032 ^ w20993;
	assign w20992 = w21022 ^ w20985;
	assign w21068 = w20989 ^ w20992;
	assign w21064 = w20985 ^ w20986;
	assign w21062 = w21072 & w21101;
	assign w21056 = w21064 & w21097;
	assign w21041 = w21056 ^ w44252;
	assign w21017 = w21056 ^ w21059;
	assign w21014 = ~w21017;
	assign w21013 = w21056 ^ w21057;
	assign w21007 = w21052 ^ w21041;
	assign w21004 = ~w21007;
	assign w21001 = w21057 ^ w21041;
	assign w21055 = w21068 & w21100;
	assign w21033 = w21051 ^ w21055;
	assign w21011 = ~w21033;
	assign w21010 = w21011 ^ w21049;
	assign w21006 = w21010 ^ w44253;
	assign w21009 = w21048 ^ w21006;
	assign w21053 = w21072 & w21103;
	assign w21047 = w21064 & w21112;
	assign w21046 = w21068 & w21109;
	assign w21012 = w21057 ^ w21046;
	assign w21008 = ~w21012;
	assign w21113 = w21008 ^ w21009;
	assign w44251 = w21047 ^ w21048;
	assign w21029 = w21053 ^ w44251;
	assign w21005 = w21029 ^ w21006;
	assign w48658 = w21004 ^ w21005;
	assign w21030 = w21054 ^ w21029;
	assign w48661 = w21030 ^ w21001;
	assign w21034 = w21062 ^ w21030;
	assign w21003 = w21061 ^ w21034;
	assign w48659 = w21002 ^ w21003;
	assign w21039 = w21063 ^ w21034;
	assign w21114 = w21039 ^ w21013;
	assign w48660 = w44252 ^ w21039;
	assign w21016 = w21020 ^ w44251;
	assign w21019 = w44253 ^ w21016;
	assign w21116 = w21018 ^ w21019;
	assign w21015 = w21011 ^ w21016;
	assign w21115 = w21014 ^ w21015;
	assign w45470 = ~w21116;
	assign w45475 = ~w21113;
	assign w45476 = ~w21114;
	assign w6560 = w48661 ^ w45476;
	assign w45477 = ~w21115;
	assign w45504 = ~w22051;
	assign w5975 = w45504 ^ w48444;
	assign w6111 = w5975 ^ w5976;
	assign w6099 = w5975 ^ w45176;
	assign w48330 = w6099 ^ w6098;
	assign w47743 = w48330 ^ w21;
	assign w45505 = ~w22052;
	assign w5977 = w45505 ^ w48445;
	assign w6101 = w5977 ^ w5533;
	assign w6086 = w5977 ^ w6028;
	assign w48324 = w48440 ^ w6086;
	assign w47749 = w48324 ^ w15;
	assign w33974 = w47752 ^ w47749;
	assign w45570 = ~w25937;
	assign w6006 = w45570 ^ w45188;
	assign w6164 = w6006 ^ w6010;
	assign w48370 = w45179 ^ w6164;
	assign w47703 = w48370 ^ w61;
	assign w45571 = ~w25938;
	assign w6139 = w48460 ^ w45571;
	assign w48356 = w6140 ^ w6139;
	assign w47717 = w48356 ^ w47;
	assign w45572 = ~w25939;
	assign w6116 = w48462 ^ w45572;
	assign w5991 = w45572 ^ w48461;
	assign w6131 = w5991 ^ w6000;
	assign w48351 = w48457 ^ w6131;
	assign w47722 = w48351 ^ w42;
	assign w35983 = w47717 ^ w47722;
	assign w45573 = ~w25940;
	assign w5990 = w45573 ^ w45190;
	assign w6275 = w5936 ^ w45573;
	assign w6151 = w5990 ^ w6031;
	assign w48365 = w45174 ^ w6151;
	assign w47708 = w48365 ^ w56;
	assign w6141 = w5990 ^ w6023;
	assign w45654 = ~w29022;
	assign w48317 = w45654 ^ w6212;
	assign w6234 = w45498 ^ w45654;
	assign w5959 = w6235 ^ w6234;
	assign w47756 = w48317 ^ w8;
	assign w45660 = ~w29019;
	assign w48338 = w45660 ^ w6111;
	assign w6100 = w45660 ^ w36121;
	assign w48331 = w6101 ^ w6100;
	assign w5980 = w45660 ^ w45176;
	assign w6084 = w5972 ^ w5980;
	assign w6157 = w5980 ^ w48439;
	assign w6159 = ~w6157;
	assign w6113 = w5977 ^ w5980;
	assign w48314 = w6159 ^ w6158;
	assign w47742 = w48331 ^ w22;
	assign w32280 = w47744 ^ w47742;
	assign w32239 = w32280 ^ w47743;
	assign w47759 = w48314 ^ w5;
	assign w47735 = w48338 ^ w29;
	assign w48322 = w45504 ^ w6084;
	assign w47751 = w48322 ^ w13;
	assign w33886 = w47751 ^ w47749;
	assign w45661 = ~w29020;
	assign w48339 = w45661 ^ w6113;
	assign w6102 = w45661 ^ w36122;
	assign w48332 = w6103 ^ w6102;
	assign w5983 = w45661 ^ w48455;
	assign w6085 = w5975 ^ w5983;
	assign w48323 = w45505 ^ w6085;
	assign w6114 = w5983 ^ w6027;
	assign w48340 = w48451 ^ w6114;
	assign w6176 = w5983 ^ w45504;
	assign w6177 = w6176 ^ w6175;
	assign w48315 = ~w6177;
	assign w47733 = w48340 ^ w31;
	assign w21290 = w47735 ^ w47733;
	assign w21377 = w47733 ^ w47738;
	assign w47750 = w48323 ^ w14;
	assign w33888 = w47752 ^ w47750;
	assign w33892 = w47756 ^ w47750;
	assign w33969 = w33886 ^ w33892;
	assign w33972 = w47751 ^ w33892;
	assign w33848 = w33888 ^ w33886;
	assign w33847 = w33888 ^ w47751;
	assign w33971 = w47756 ^ w33847;
	assign w33957 = w47756 & w33971;
	assign w47741 = w48332 ^ w23;
	assign w32278 = w47743 ^ w47741;
	assign w32366 = w47744 ^ w47741;
	assign w32240 = w32280 ^ w32278;
	assign w47734 = w48339 ^ w30;
	assign w47758 = w48315 ^ w6;
	assign w32414 = w47760 ^ w47758;
	assign w32373 = w32414 ^ w47759;
	assign w45754 = ~w32640;
	assign w5993 = w45174 ^ w45754;
	assign w6127 = w5993 ^ w6030;
	assign w48349 = w45573 ^ w6127;
	assign w6115 = w5993 ^ w6021;
	assign w48341 = w45190 ^ w6115;
	assign w6153 = w5991 ^ w5993;
	assign w6276 = w6274 ^ w45754;
	assign w5942 = w6276 ^ w6275;
	assign w47724 = w48349 ^ w40;
	assign w47732 = w48341 ^ w32;
	assign w48357 = w45754 ^ w6141;
	assign w47716 = w48357 ^ w48;
	assign w48366 = w6153 ^ w6152;
	assign w47707 = w48366 ^ w57;
	assign w25711 = w47707 ^ w47705;
	assign w45759 = ~w32637;
	assign w6145 = w6006 ^ w45759;
	assign w6147 = ~w6145;
	assign w6120 = w45759 ^ w45570;
	assign w48362 = w6147 ^ w6146;
	assign w47711 = w48362 ^ w53;
	assign w21156 = w47711 ^ w47709;
	assign w21231 = w21156 ^ w21246;
	assign w21222 = w21246 & w21231;
	assign w6015 = w45179 ^ w45759;
	assign w6119 = w6015 ^ w48472;
	assign w48346 = w6119 ^ w6118;
	assign w6137 = w6002 ^ w6015;
	assign w48354 = w45570 ^ w6137;
	assign w47719 = w48354 ^ w45;
	assign w35896 = w47719 ^ w47717;
	assign w47727 = w48346 ^ w37;
	assign w6165 = w6013 ^ w6015;
	assign w48371 = w45571 ^ w6165;
	assign w47702 = w48371 ^ w62;
	assign w25714 = w47704 ^ w47702;
	assign w25718 = w47708 ^ w47702;
	assign w25798 = w47703 ^ w25718;
	assign w25794 = w47707 ^ w25798;
	assign w25673 = w25714 ^ w47703;
	assign w25797 = w47708 ^ w25673;
	assign w25783 = w47708 & w25797;
	assign w25781 = w25798 & w25794;
	assign w45760 = ~w32638;
	assign w6121 = w6013 ^ w45760;
	assign w6167 = w6030 ^ w45760;
	assign w48372 = w6167 ^ w6166;
	assign w48347 = w6121 ^ w6120;
	assign w47701 = w48372 ^ w63;
	assign w6012 = w45571 ^ w45760;
	assign w6122 = w6012 ^ w6031;
	assign w48348 = w48465 ^ w6122;
	assign w6149 = w6012 ^ w45179;
	assign w25712 = w47703 ^ w47701;
	assign w25800 = w47704 ^ w47701;
	assign w25795 = w25712 ^ w25718;
	assign w25792 = w25711 ^ w25800;
	assign w25791 = w47708 ^ w25792;
	assign w25674 = w25714 ^ w25712;
	assign w25790 = w25711 ^ w25674;
	assign w25801 = w47701 ^ w47707;
	assign w48363 = w6149 ^ w6148;
	assign w6138 = w6006 ^ w6012;
	assign w47710 = w48363 ^ w54;
	assign w21158 = w47712 ^ w47710;
	assign w21162 = w47716 ^ w47710;
	assign w21239 = w21156 ^ w21162;
	assign w21242 = w47711 ^ w21162;
	assign w21118 = w21158 ^ w21156;
	assign w21117 = w21158 ^ w47711;
	assign w21241 = w47716 ^ w21117;
	assign w21227 = w47716 & w21241;
	assign w47726 = w48347 ^ w38;
	assign w28796 = w47728 ^ w47726;
	assign w28800 = w47732 ^ w47726;
	assign w28880 = w47727 ^ w28800;
	assign w28755 = w28796 ^ w47727;
	assign w28879 = w47732 ^ w28755;
	assign w28865 = w47732 & w28879;
	assign w47725 = w48348 ^ w39;
	assign w28794 = w47727 ^ w47725;
	assign w28882 = w47728 ^ w47725;
	assign w28877 = w28794 ^ w28800;
	assign w28756 = w28796 ^ w28794;
	assign w48355 = w45172 ^ w6138;
	assign w47718 = w48355 ^ w46;
	assign w35902 = w47724 ^ w47718;
	assign w35979 = w35896 ^ w35902;
	assign w35982 = w47719 ^ w35902;
	assign w45761 = ~w32639;
	assign w6117 = w6000 ^ w45761;
	assign w48343 = w6117 ^ w6116;
	assign w5997 = w45173 ^ w45761;
	assign w6129 = w5990 ^ w5997;
	assign w48342 = w5942 ^ w5997;
	assign w6154 = w5995 ^ w5997;
	assign w6264 = w6023 ^ w45761;
	assign w5947 = w6264 ^ w6263;
	assign w48358 = w5947 ^ w5991;
	assign w47715 = w48358 ^ w49;
	assign w21155 = w47715 ^ w47713;
	assign w21157 = w47714 ^ w21155;
	assign w21233 = w47710 ^ w21157;
	assign w21230 = w47711 ^ w21157;
	assign w21232 = w21162 ^ w21157;
	assign w21238 = w47715 ^ w21242;
	assign w21236 = w21155 ^ w21244;
	assign w21235 = w47716 ^ w21236;
	assign w21172 = w47715 ^ w47714;
	assign w21237 = w21172 ^ w21239;
	assign w21240 = w21244 ^ w21172;
	assign w21234 = w21155 ^ w21118;
	assign w21245 = w47709 ^ w47715;
	assign w21229 = w21236 & w21240;
	assign w21161 = w21229 ^ w21158;
	assign w21228 = w21237 & w21235;
	assign w21179 = w21222 ^ w21228;
	assign w21226 = w21245 & w21230;
	assign w21160 = w21226 ^ w21156;
	assign w21225 = w21242 & w21238;
	assign w21224 = w21239 & w21232;
	assign w21223 = w21244 & w21233;
	assign w21159 = w21223 ^ w21157;
	assign w21165 = w21161 ^ w21159;
	assign w21170 = w47709 ^ w21165;
	assign w21220 = w21179 ^ w21170;
	assign w21131 = w21222 ^ w21223;
	assign w21178 = w21131 ^ w21132;
	assign w21177 = w21178 ^ w21160;
	assign w21219 = w21225 ^ w21177;
	assign w21221 = w21243 & w21234;
	assign w21216 = w21220 & w21219;
	assign w47731 = w48342 ^ w33;
	assign w28793 = w47731 ^ w47729;
	assign w28876 = w47731 ^ w28880;
	assign w28874 = w28793 ^ w28882;
	assign w28873 = w47732 ^ w28874;
	assign w28872 = w28793 ^ w28756;
	assign w28883 = w47725 ^ w47731;
	assign w28863 = w28880 & w28876;
	assign w47730 = w48343 ^ w34;
	assign w28795 = w47730 ^ w28793;
	assign w28871 = w47726 ^ w28795;
	assign w28868 = w47727 ^ w28795;
	assign w28870 = w28800 ^ w28795;
	assign w28810 = w47731 ^ w47730;
	assign w28875 = w28810 ^ w28877;
	assign w28878 = w28882 ^ w28810;
	assign w28884 = w47730 ^ w47728;
	assign w28869 = w28794 ^ w28884;
	assign w28770 = w47729 ^ w47730;
	assign w28881 = w47725 ^ w47730;
	assign w28867 = w28874 & w28878;
	assign w28799 = w28867 ^ w28796;
	assign w28866 = w28875 & w28873;
	assign w28864 = w28883 & w28868;
	assign w28798 = w28864 ^ w28794;
	assign w28862 = w28877 & w28870;
	assign w28861 = w28882 & w28871;
	assign w28797 = w28861 ^ w28795;
	assign w28803 = w28799 ^ w28797;
	assign w28808 = w47725 ^ w28803;
	assign w28860 = w28884 & w28869;
	assign w28817 = w28860 ^ w28866;
	assign w28858 = w28817 ^ w28808;
	assign w28769 = w28860 ^ w28861;
	assign w28816 = w28769 ^ w28770;
	assign w28815 = w28816 ^ w28798;
	assign w28857 = w28863 ^ w28815;
	assign w28859 = w28881 & w28872;
	assign w28854 = w28858 & w28857;
	assign w44255 = w21221 ^ w21224;
	assign w21134 = w21160 ^ w44255;
	assign w21218 = w21134 ^ w21159;
	assign w21215 = w21216 ^ w21218;
	assign w21174 = w21222 ^ w44255;
	assign w21130 = w21225 ^ w21174;
	assign w21212 = w47715 ^ w21130;
	assign w44258 = w21221 ^ w21227;
	assign w21133 = w21165 ^ w44258;
	assign w21176 = w47711 ^ w21133;
	assign w21211 = w21216 ^ w21176;
	assign w21210 = w21211 & w21212;
	assign w21209 = w21210 ^ w21218;
	assign w21208 = w21216 ^ w21210;
	assign w21129 = w21210 ^ w21174;
	assign w21128 = w21210 ^ w21227;
	assign w21123 = w21128 ^ w21224;
	assign w21207 = w21218 & w21208;
	assign w21205 = w21207 ^ w21215;
	assign w21195 = w21209 & w47716;
	assign w21186 = w21209 & w21241;
	assign w44257 = w21207 ^ w21225;
	assign w21199 = w44257 ^ w21177;
	assign w21197 = w21199 & w21236;
	assign w21188 = w21199 & w21240;
	assign w21166 = w47715 ^ w44257;
	assign w21206 = w21166 ^ w21129;
	assign w21196 = w21206 & w21235;
	assign w21187 = w21206 & w21237;
	assign w21171 = w44258 ^ w21156;
	assign w21217 = w21179 ^ w21171;
	assign w21214 = w21217 & w21215;
	assign w21213 = w21214 ^ w21176;
	assign w21125 = w21214 ^ w21226;
	assign w21121 = w21125 ^ w21161;
	assign w21124 = w47709 ^ w21121;
	assign w21201 = w21123 ^ w21124;
	assign w21122 = w21214 ^ w21170;
	assign w21120 = w47711 ^ w21121;
	assign w21204 = w21213 & w21205;
	assign w21169 = w21204 ^ w21179;
	assign w21203 = w21169 ^ w21171;
	assign w21127 = w21204 ^ w21228;
	assign w21119 = w21166 ^ w21127;
	assign w21126 = w21156 ^ w21119;
	assign w21202 = w21123 ^ w21126;
	assign w21200 = w21169 ^ w21122;
	assign w21198 = w21119 ^ w21120;
	assign w21194 = w21200 & w21230;
	assign w21193 = w21203 & w21242;
	assign w21192 = w21213 & w21232;
	assign w21136 = w21192 ^ w21193;
	assign w21191 = w21201 & w21233;
	assign w21190 = w21198 & w21231;
	assign w21151 = w21190 ^ w21193;
	assign w21148 = ~w21151;
	assign w21147 = w21190 ^ w21191;
	assign w21189 = w21202 & w21234;
	assign w21185 = w21200 & w21245;
	assign w21167 = w21185 ^ w21189;
	assign w21152 = w21194 ^ w21185;
	assign w21145 = ~w21167;
	assign w21184 = w21203 & w21238;
	assign w21154 = w21192 ^ w21184;
	assign w21183 = w21213 & w21239;
	assign w21144 = w21145 ^ w21183;
	assign w21182 = w21201 & w21244;
	assign w21181 = w21198 & w21246;
	assign w21180 = w21202 & w21243;
	assign w21146 = w21191 ^ w21180;
	assign w21142 = ~w21146;
	assign w44256 = w21181 ^ w21182;
	assign w21163 = w21187 ^ w44256;
	assign w21164 = w21188 ^ w21163;
	assign w21168 = w21196 ^ w21164;
	assign w21173 = w21197 ^ w21168;
	assign w21248 = w21173 ^ w21147;
	assign w21137 = w21195 ^ w21168;
	assign w48687 = w21136 ^ w21137;
	assign w21150 = w21154 ^ w44256;
	assign w21149 = w21145 ^ w21150;
	assign w21249 = w21148 ^ w21149;
	assign w44259 = w21193 ^ w21194;
	assign w48688 = w44259 ^ w21173;
	assign w21175 = w21190 ^ w44259;
	assign w21141 = w21186 ^ w21175;
	assign w21138 = ~w21141;
	assign w21135 = w21191 ^ w21175;
	assign w48689 = w21164 ^ w21135;
	assign w44260 = w21195 ^ w21197;
	assign w21153 = w44260 ^ w21150;
	assign w21250 = w21152 ^ w21153;
	assign w21140 = w21144 ^ w44260;
	assign w21143 = w21182 ^ w21140;
	assign w21247 = w21142 ^ w21143;
	assign w21139 = w21163 ^ w21140;
	assign w48686 = w21138 ^ w21139;
	assign w48367 = w48466 ^ w6154;
	assign w47706 = w48367 ^ w58;
	assign w25713 = w47706 ^ w25711;
	assign w25789 = w47702 ^ w25713;
	assign w25786 = w47703 ^ w25713;
	assign w25788 = w25718 ^ w25713;
	assign w25728 = w47707 ^ w47706;
	assign w25793 = w25728 ^ w25795;
	assign w25796 = w25800 ^ w25728;
	assign w25802 = w47706 ^ w47704;
	assign w25787 = w25712 ^ w25802;
	assign w25688 = w47705 ^ w47706;
	assign w25799 = w47701 ^ w47706;
	assign w25785 = w25792 & w25796;
	assign w25717 = w25785 ^ w25714;
	assign w25784 = w25793 & w25791;
	assign w25782 = w25801 & w25786;
	assign w25716 = w25782 ^ w25712;
	assign w25780 = w25795 & w25788;
	assign w25779 = w25800 & w25789;
	assign w25715 = w25779 ^ w25713;
	assign w25721 = w25717 ^ w25715;
	assign w25726 = w47701 ^ w25721;
	assign w25778 = w25802 & w25787;
	assign w25735 = w25778 ^ w25784;
	assign w25776 = w25735 ^ w25726;
	assign w25687 = w25778 ^ w25779;
	assign w25734 = w25687 ^ w25688;
	assign w25733 = w25734 ^ w25716;
	assign w25775 = w25781 ^ w25733;
	assign w25777 = w25799 & w25790;
	assign w25772 = w25776 & w25775;
	assign w44446 = w25777 ^ w25780;
	assign w25690 = w25716 ^ w44446;
	assign w25774 = w25690 ^ w25715;
	assign w25771 = w25772 ^ w25774;
	assign w25730 = w25778 ^ w44446;
	assign w25686 = w25781 ^ w25730;
	assign w25768 = w47707 ^ w25686;
	assign w44449 = w25777 ^ w25783;
	assign w25689 = w25721 ^ w44449;
	assign w25732 = w47703 ^ w25689;
	assign w25767 = w25772 ^ w25732;
	assign w25766 = w25767 & w25768;
	assign w25765 = w25766 ^ w25774;
	assign w25764 = w25772 ^ w25766;
	assign w25685 = w25766 ^ w25730;
	assign w25684 = w25766 ^ w25783;
	assign w25679 = w25684 ^ w25780;
	assign w25763 = w25774 & w25764;
	assign w25761 = w25763 ^ w25771;
	assign w25751 = w25765 & w47708;
	assign w25742 = w25765 & w25797;
	assign w44448 = w25763 ^ w25781;
	assign w25755 = w44448 ^ w25733;
	assign w25753 = w25755 & w25792;
	assign w25744 = w25755 & w25796;
	assign w25722 = w47707 ^ w44448;
	assign w25762 = w25722 ^ w25685;
	assign w25752 = w25762 & w25791;
	assign w25743 = w25762 & w25793;
	assign w25727 = w44449 ^ w25712;
	assign w25773 = w25735 ^ w25727;
	assign w25770 = w25773 & w25771;
	assign w25769 = w25770 ^ w25732;
	assign w25681 = w25770 ^ w25782;
	assign w25677 = w25681 ^ w25717;
	assign w25680 = w47701 ^ w25677;
	assign w25757 = w25679 ^ w25680;
	assign w25678 = w25770 ^ w25726;
	assign w25676 = w47703 ^ w25677;
	assign w25760 = w25769 & w25761;
	assign w25725 = w25760 ^ w25735;
	assign w25759 = w25725 ^ w25727;
	assign w25683 = w25760 ^ w25784;
	assign w25675 = w25722 ^ w25683;
	assign w25682 = w25712 ^ w25675;
	assign w25758 = w25679 ^ w25682;
	assign w25756 = w25725 ^ w25678;
	assign w25754 = w25675 ^ w25676;
	assign w25750 = w25756 & w25786;
	assign w25749 = w25759 & w25798;
	assign w25748 = w25769 & w25788;
	assign w25692 = w25748 ^ w25749;
	assign w25747 = w25757 & w25789;
	assign w25746 = w25754 & w25787;
	assign w25707 = w25746 ^ w25749;
	assign w25704 = ~w25707;
	assign w25703 = w25746 ^ w25747;
	assign w25745 = w25758 & w25790;
	assign w25741 = w25756 & w25801;
	assign w25723 = w25741 ^ w25745;
	assign w25708 = w25750 ^ w25741;
	assign w25701 = ~w25723;
	assign w25740 = w25759 & w25794;
	assign w25710 = w25748 ^ w25740;
	assign w25739 = w25769 & w25795;
	assign w25700 = w25701 ^ w25739;
	assign w25738 = w25757 & w25800;
	assign w25737 = w25754 & w25802;
	assign w25736 = w25758 & w25799;
	assign w25702 = w25747 ^ w25736;
	assign w25698 = ~w25702;
	assign w44447 = w25737 ^ w25738;
	assign w25719 = w25743 ^ w44447;
	assign w25720 = w25744 ^ w25719;
	assign w25724 = w25752 ^ w25720;
	assign w25729 = w25753 ^ w25724;
	assign w25804 = w25729 ^ w25703;
	assign w25693 = w25751 ^ w25724;
	assign w48672 = w25692 ^ w25693;
	assign w25706 = w25710 ^ w44447;
	assign w25705 = w25701 ^ w25706;
	assign w25805 = w25704 ^ w25705;
	assign w44450 = w25749 ^ w25750;
	assign w48673 = w44450 ^ w25729;
	assign w25731 = w25746 ^ w44450;
	assign w25697 = w25742 ^ w25731;
	assign w25694 = ~w25697;
	assign w25691 = w25747 ^ w25731;
	assign w48674 = w25720 ^ w25691;
	assign w6678 = w48661 ^ w48674;
	assign w6429 = w6678 ^ w48672;
	assign w6425 = ~w6678;
	assign w44451 = w25751 ^ w25753;
	assign w25709 = w44451 ^ w25706;
	assign w25806 = w25708 ^ w25709;
	assign w25696 = w25700 ^ w44451;
	assign w25699 = w25738 ^ w25696;
	assign w25803 = w25698 ^ w25699;
	assign w25695 = w25719 ^ w25696;
	assign w48671 = w25694 ^ w25695;
	assign w6426 = w6425 ^ w48671;
	assign w44574 = w28859 ^ w28865;
	assign w28771 = w28803 ^ w44574;
	assign w28814 = w47727 ^ w28771;
	assign w28849 = w28854 ^ w28814;
	assign w28809 = w44574 ^ w28794;
	assign w28855 = w28817 ^ w28809;
	assign w44575 = w28859 ^ w28862;
	assign w28812 = w28860 ^ w44575;
	assign w28768 = w28863 ^ w28812;
	assign w28850 = w47731 ^ w28768;
	assign w28848 = w28849 & w28850;
	assign w28766 = w28848 ^ w28865;
	assign w28767 = w28848 ^ w28812;
	assign w28846 = w28854 ^ w28848;
	assign w28761 = w28766 ^ w28862;
	assign w28772 = w28798 ^ w44575;
	assign w28856 = w28772 ^ w28797;
	assign w28847 = w28848 ^ w28856;
	assign w28853 = w28854 ^ w28856;
	assign w28852 = w28855 & w28853;
	assign w28851 = w28852 ^ w28814;
	assign w28763 = w28852 ^ w28864;
	assign w28759 = w28763 ^ w28799;
	assign w28762 = w47725 ^ w28759;
	assign w28839 = w28761 ^ w28762;
	assign w28760 = w28852 ^ w28808;
	assign w28758 = w47727 ^ w28759;
	assign w28845 = w28856 & w28846;
	assign w28843 = w28845 ^ w28853;
	assign w28842 = w28851 & w28843;
	assign w28807 = w28842 ^ w28817;
	assign w28841 = w28807 ^ w28809;
	assign w28765 = w28842 ^ w28866;
	assign w28838 = w28807 ^ w28760;
	assign w28833 = w28847 & w47732;
	assign w28832 = w28838 & w28868;
	assign w28831 = w28841 & w28880;
	assign w28830 = w28851 & w28870;
	assign w28774 = w28830 ^ w28831;
	assign w28829 = w28839 & w28871;
	assign w28824 = w28847 & w28879;
	assign w28823 = w28838 & w28883;
	assign w28790 = w28832 ^ w28823;
	assign w28822 = w28841 & w28876;
	assign w28792 = w28830 ^ w28822;
	assign w28821 = w28851 & w28877;
	assign w28820 = w28839 & w28882;
	assign w44577 = w28831 ^ w28832;
	assign w44579 = w28845 ^ w28863;
	assign w28837 = w44579 ^ w28815;
	assign w28835 = w28837 & w28874;
	assign w44578 = w28833 ^ w28835;
	assign w28826 = w28837 & w28878;
	assign w28804 = w47731 ^ w44579;
	assign w28844 = w28804 ^ w28767;
	assign w28757 = w28804 ^ w28765;
	assign w28764 = w28794 ^ w28757;
	assign w28840 = w28761 ^ w28764;
	assign w28836 = w28757 ^ w28758;
	assign w28834 = w28844 & w28873;
	assign w28828 = w28836 & w28869;
	assign w28813 = w28828 ^ w44577;
	assign w28789 = w28828 ^ w28831;
	assign w28786 = ~w28789;
	assign w28785 = w28828 ^ w28829;
	assign w28779 = w28824 ^ w28813;
	assign w28776 = ~w28779;
	assign w28773 = w28829 ^ w28813;
	assign w28827 = w28840 & w28872;
	assign w28805 = w28823 ^ w28827;
	assign w28783 = ~w28805;
	assign w28782 = w28783 ^ w28821;
	assign w28778 = w28782 ^ w44578;
	assign w28781 = w28820 ^ w28778;
	assign w28825 = w28844 & w28875;
	assign w28819 = w28836 & w28884;
	assign w28818 = w28840 & w28881;
	assign w28784 = w28829 ^ w28818;
	assign w28780 = ~w28784;
	assign w28885 = w28780 ^ w28781;
	assign w44576 = w28819 ^ w28820;
	assign w28801 = w28825 ^ w44576;
	assign w28777 = w28801 ^ w28778;
	assign w48638 = w28776 ^ w28777;
	assign w28802 = w28826 ^ w28801;
	assign w48641 = w28802 ^ w28773;
	assign w28806 = w28834 ^ w28802;
	assign w28775 = w28833 ^ w28806;
	assign w48639 = w28774 ^ w28775;
	assign w28811 = w28835 ^ w28806;
	assign w28886 = w28811 ^ w28785;
	assign w48640 = w44577 ^ w28811;
	assign w28788 = w28792 ^ w44576;
	assign w28791 = w44578 ^ w28788;
	assign w28888 = w28790 ^ w28791;
	assign w28787 = w28783 ^ w28788;
	assign w28887 = w28786 ^ w28787;
	assign w45474 = ~w21250;
	assign w45479 = ~w21247;
	assign w45480 = ~w21248;
	assign w45481 = ~w21249;
	assign w45566 = ~w25803;
	assign w6579 = w45566 ^ w45475;
	assign w45567 = ~w25804;
	assign w6687 = w45476 ^ w45567;
	assign w45568 = ~w25805;
	assign w45569 = ~w25806;
	assign w6423 = w6425 ^ w45569;
	assign w45650 = ~w28888;
	assign w45655 = ~w28885;
	assign w45656 = ~w28886;
	assign w45657 = ~w28887;
	assign w45798 = ~w38670;
	assign w48413 = w45798 ^ w6044;
	assign w5971 = w45798 ^ w45183;
	assign w6059 = w5971 ^ w6019;
	assign w48421 = w45483 ^ w6059;
	assign w6069 = w5971 ^ w6034;
	assign w48429 = w45491 ^ w6069;
	assign w6046 = w5971 ^ w6004;
	assign w6268 = w6022 ^ w45798;
	assign w5945 = w6268 ^ w6267;
	assign w48406 = w5945 ^ w6004;
	assign w47667 = w48406 ^ w97;
	assign w20887 = w47667 ^ w47665;
	assign w47660 = w48413 ^ w104;
	assign w47652 = w48421 ^ w112;
	assign w20760 = w47652 ^ w47646;
	assign w47644 = w48429 ^ w120;
	assign w32016 = w47644 ^ w47638;
	assign w45799 = ~w36123;
	assign w6054 = w6123 ^ w45799;
	assign w6088 = w6092 ^ w45799;
	assign w48319 = w6054 ^ w6053;
	assign w5986 = w45799 ^ w48447;
	assign w6091 = w5985 ^ w5986;
	assign w48327 = w48441 ^ w6091;
	assign w6096 = w5964 ^ w5986;
	assign w6097 = w6096 ^ w6095;
	assign w48310 = ~w6097;
	assign w48334 = w5959 ^ w5986;
	assign w47754 = w48319 ^ w10;
	assign w33976 = w47754 ^ w47752;
	assign w33961 = w33886 ^ w33976;
	assign w33862 = w47753 ^ w47754;
	assign w33973 = w47749 ^ w47754;
	assign w33952 = w33976 & w33961;
	assign w47746 = w48327 ^ w18;
	assign w32368 = w47746 ^ w47744;
	assign w32353 = w32278 ^ w32368;
	assign w32254 = w47745 ^ w47746;
	assign w32365 = w47741 ^ w47746;
	assign w32344 = w32368 & w32353;
	assign w47739 = w48334 ^ w25;
	assign w21306 = w47739 ^ w47738;
	assign w21379 = w47733 ^ w47739;
	assign w47763 = w48310 ^ w1;
	assign w32411 = w47763 ^ w47761;
	assign w32413 = w47762 ^ w32411;
	assign w32489 = w47758 ^ w32413;
	assign w32486 = w47759 ^ w32413;
	assign w32428 = w47763 ^ w47762;
	assign w45800 = ~w36124;
	assign w48325 = w45800 ^ w6087;
	assign w5987 = w45800 ^ w45654;
	assign w6089 = w5965 ^ w5987;
	assign w6104 = w5987 ^ w6028;
	assign w48333 = w45499 ^ w6104;
	assign w6090 = w6089 ^ w6088;
	assign w48326 = ~w6090;
	assign w6035 = w5987 ^ w6020;
	assign w48309 = w45178 ^ w6035;
	assign w6239 = w5938 ^ w45800;
	assign w47747 = w48326 ^ w17;
	assign w32277 = w47747 ^ w47745;
	assign w32279 = w47746 ^ w32277;
	assign w32355 = w47742 ^ w32279;
	assign w32352 = w47743 ^ w32279;
	assign w32358 = w32277 ^ w32366;
	assign w32294 = w47747 ^ w47746;
	assign w32362 = w32366 ^ w32294;
	assign w32356 = w32277 ^ w32240;
	assign w32367 = w47741 ^ w47747;
	assign w32351 = w32358 & w32362;
	assign w32283 = w32351 ^ w32280;
	assign w32348 = w32367 & w32352;
	assign w32282 = w32348 ^ w32278;
	assign w32345 = w32366 & w32355;
	assign w32281 = w32345 ^ w32279;
	assign w32287 = w32283 ^ w32281;
	assign w32292 = w47741 ^ w32287;
	assign w32253 = w32344 ^ w32345;
	assign w32300 = w32253 ^ w32254;
	assign w32299 = w32300 ^ w32282;
	assign w32343 = w32365 & w32356;
	assign w47764 = w48309 ^ w0;
	assign w32418 = w47764 ^ w47758;
	assign w32488 = w32418 ^ w32413;
	assign w32498 = w47759 ^ w32418;
	assign w32494 = w47763 ^ w32498;
	assign w32497 = w47764 ^ w32373;
	assign w32483 = w47764 & w32497;
	assign w32481 = w32498 & w32494;
	assign w47740 = w48333 ^ w24;
	assign w21296 = w47740 ^ w47734;
	assign w21373 = w21290 ^ w21296;
	assign w21371 = w21306 ^ w21373;
	assign w21376 = w47735 ^ w21296;
	assign w21372 = w47739 ^ w21376;
	assign w21359 = w21376 & w21372;
	assign w47748 = w48325 ^ w16;
	assign w32357 = w47748 ^ w32358;
	assign w32284 = w47748 ^ w47742;
	assign w32354 = w32284 ^ w32279;
	assign w32361 = w32278 ^ w32284;
	assign w32359 = w32294 ^ w32361;
	assign w32364 = w47743 ^ w32284;
	assign w32360 = w47747 ^ w32364;
	assign w32363 = w47748 ^ w32239;
	assign w32350 = w32359 & w32357;
	assign w32301 = w32344 ^ w32350;
	assign w32342 = w32301 ^ w32292;
	assign w32349 = w47748 & w32363;
	assign w32347 = w32364 & w32360;
	assign w32341 = w32347 ^ w32299;
	assign w32346 = w32361 & w32354;
	assign w32338 = w32342 & w32341;
	assign w44722 = w32343 ^ w32349;
	assign w32293 = w44722 ^ w32278;
	assign w32339 = w32301 ^ w32293;
	assign w32255 = w32287 ^ w44722;
	assign w32298 = w47743 ^ w32255;
	assign w32333 = w32338 ^ w32298;
	assign w44723 = w32343 ^ w32346;
	assign w32296 = w32344 ^ w44723;
	assign w32252 = w32347 ^ w32296;
	assign w32334 = w47747 ^ w32252;
	assign w32332 = w32333 & w32334;
	assign w32251 = w32332 ^ w32296;
	assign w32250 = w32332 ^ w32349;
	assign w32245 = w32250 ^ w32346;
	assign w32330 = w32338 ^ w32332;
	assign w32256 = w32282 ^ w44723;
	assign w32340 = w32256 ^ w32281;
	assign w32331 = w32332 ^ w32340;
	assign w32337 = w32338 ^ w32340;
	assign w32336 = w32339 & w32337;
	assign w32335 = w32336 ^ w32298;
	assign w32247 = w32336 ^ w32348;
	assign w32243 = w32247 ^ w32283;
	assign w32246 = w47741 ^ w32243;
	assign w32323 = w32245 ^ w32246;
	assign w32244 = w32336 ^ w32292;
	assign w32242 = w47743 ^ w32243;
	assign w32329 = w32340 & w32330;
	assign w32327 = w32329 ^ w32337;
	assign w32326 = w32335 & w32327;
	assign w32291 = w32326 ^ w32301;
	assign w32325 = w32291 ^ w32293;
	assign w32249 = w32326 ^ w32350;
	assign w32322 = w32291 ^ w32244;
	assign w32317 = w32331 & w47748;
	assign w32316 = w32322 & w32352;
	assign w32315 = w32325 & w32364;
	assign w32314 = w32335 & w32354;
	assign w32258 = w32314 ^ w32315;
	assign w32313 = w32323 & w32355;
	assign w32308 = w32331 & w32363;
	assign w32307 = w32322 & w32367;
	assign w32274 = w32316 ^ w32307;
	assign w32306 = w32325 & w32360;
	assign w32276 = w32314 ^ w32306;
	assign w32305 = w32335 & w32361;
	assign w32304 = w32323 & w32366;
	assign w44724 = w32315 ^ w32316;
	assign w44726 = w32329 ^ w32347;
	assign w32288 = w47747 ^ w44726;
	assign w32328 = w32288 ^ w32251;
	assign w32309 = w32328 & w32359;
	assign w32318 = w32328 & w32357;
	assign w32241 = w32288 ^ w32249;
	assign w32248 = w32278 ^ w32241;
	assign w32324 = w32245 ^ w32248;
	assign w32311 = w32324 & w32356;
	assign w32289 = w32307 ^ w32311;
	assign w32267 = ~w32289;
	assign w32266 = w32267 ^ w32305;
	assign w32320 = w32241 ^ w32242;
	assign w32303 = w32320 & w32368;
	assign w32302 = w32324 & w32365;
	assign w32268 = w32313 ^ w32302;
	assign w32264 = ~w32268;
	assign w43589 = w32303 ^ w32304;
	assign w32272 = w32276 ^ w43589;
	assign w32271 = w32267 ^ w32272;
	assign w32285 = w32309 ^ w43589;
	assign w32312 = w32320 & w32353;
	assign w32269 = w32312 ^ w32313;
	assign w32273 = w32312 ^ w32315;
	assign w32270 = ~w32273;
	assign w32371 = w32270 ^ w32271;
	assign w32297 = w32312 ^ w44724;
	assign w32263 = w32308 ^ w32297;
	assign w32257 = w32313 ^ w32297;
	assign w32260 = ~w32263;
	assign w32321 = w44726 ^ w32299;
	assign w32319 = w32321 & w32358;
	assign w32310 = w32321 & w32362;
	assign w32286 = w32310 ^ w32285;
	assign w32290 = w32318 ^ w32286;
	assign w32295 = w32319 ^ w32290;
	assign w48669 = w44724 ^ w32295;
	assign w32370 = w32295 ^ w32269;
	assign w32259 = w32317 ^ w32290;
	assign w48668 = w32258 ^ w32259;
	assign w48670 = w32286 ^ w32257;
	assign w6689 = w48669 ^ w48673;
	assign w6538 = ~w48669;
	assign w6694 = w48668 ^ w48672;
	assign w44725 = w32317 ^ w32319;
	assign w32275 = w44725 ^ w32272;
	assign w32372 = w32274 ^ w32275;
	assign w32262 = w32266 ^ w44725;
	assign w32265 = w32304 ^ w32262;
	assign w32369 = w32264 ^ w32265;
	assign w32261 = w32285 ^ w32262;
	assign w48667 = w32260 ^ w32261;
	assign w6699 = w48667 ^ w48671;
	assign w6582 = w6699 ^ w45568;
	assign w6668 = w48670 ^ w48674;
	assign w6537 = w6668 ^ w6538;
	assign w6577 = w6687 ^ w6668;
	assign w6544 = w6668 ^ w48668;
	assign w5957 = w6239 ^ w6238;
	assign w48318 = w5957 ^ w5965;
	assign w47755 = w48318 ^ w9;
	assign w33885 = w47755 ^ w47753;
	assign w33887 = w47754 ^ w33885;
	assign w33963 = w47750 ^ w33887;
	assign w33960 = w47751 ^ w33887;
	assign w33962 = w33892 ^ w33887;
	assign w33968 = w47755 ^ w33972;
	assign w33966 = w33885 ^ w33974;
	assign w33965 = w47756 ^ w33966;
	assign w33902 = w47755 ^ w47754;
	assign w33967 = w33902 ^ w33969;
	assign w33970 = w33974 ^ w33902;
	assign w33964 = w33885 ^ w33848;
	assign w33975 = w47749 ^ w47755;
	assign w33959 = w33966 & w33970;
	assign w33891 = w33959 ^ w33888;
	assign w33958 = w33967 & w33965;
	assign w33909 = w33952 ^ w33958;
	assign w33956 = w33975 & w33960;
	assign w33890 = w33956 ^ w33886;
	assign w33955 = w33972 & w33968;
	assign w33954 = w33969 & w33962;
	assign w33953 = w33974 & w33963;
	assign w33889 = w33953 ^ w33887;
	assign w33895 = w33891 ^ w33889;
	assign w33900 = w47749 ^ w33895;
	assign w33950 = w33909 ^ w33900;
	assign w33861 = w33952 ^ w33953;
	assign w33908 = w33861 ^ w33862;
	assign w33907 = w33908 ^ w33890;
	assign w33949 = w33955 ^ w33907;
	assign w33951 = w33973 & w33964;
	assign w33946 = w33950 & w33949;
	assign w44788 = w33951 ^ w33957;
	assign w33863 = w33895 ^ w44788;
	assign w33906 = w47751 ^ w33863;
	assign w33941 = w33946 ^ w33906;
	assign w33901 = w44788 ^ w33886;
	assign w33947 = w33909 ^ w33901;
	assign w44789 = w33951 ^ w33954;
	assign w33904 = w33952 ^ w44789;
	assign w33860 = w33955 ^ w33904;
	assign w33942 = w47755 ^ w33860;
	assign w33940 = w33941 & w33942;
	assign w33859 = w33940 ^ w33904;
	assign w33938 = w33946 ^ w33940;
	assign w33858 = w33940 ^ w33957;
	assign w33853 = w33858 ^ w33954;
	assign w33864 = w33890 ^ w44789;
	assign w33948 = w33864 ^ w33889;
	assign w33939 = w33940 ^ w33948;
	assign w33945 = w33946 ^ w33948;
	assign w33944 = w33947 & w33945;
	assign w33943 = w33944 ^ w33906;
	assign w33855 = w33944 ^ w33956;
	assign w33851 = w33855 ^ w33891;
	assign w33854 = w47749 ^ w33851;
	assign w33931 = w33853 ^ w33854;
	assign w33852 = w33944 ^ w33900;
	assign w33850 = w47751 ^ w33851;
	assign w33937 = w33948 & w33938;
	assign w33935 = w33937 ^ w33945;
	assign w33934 = w33943 & w33935;
	assign w33899 = w33934 ^ w33909;
	assign w33933 = w33899 ^ w33901;
	assign w33857 = w33934 ^ w33958;
	assign w33930 = w33899 ^ w33852;
	assign w33925 = w33939 & w47756;
	assign w33924 = w33930 & w33960;
	assign w33923 = w33933 & w33972;
	assign w33922 = w33943 & w33962;
	assign w33866 = w33922 ^ w33923;
	assign w33921 = w33931 & w33963;
	assign w33916 = w33939 & w33971;
	assign w33915 = w33930 & w33975;
	assign w33882 = w33924 ^ w33915;
	assign w33914 = w33933 & w33968;
	assign w33884 = w33922 ^ w33914;
	assign w33913 = w33943 & w33969;
	assign w33912 = w33931 & w33974;
	assign w44791 = w33923 ^ w33924;
	assign w44793 = w33937 ^ w33955;
	assign w33929 = w44793 ^ w33907;
	assign w33927 = w33929 & w33966;
	assign w44792 = w33925 ^ w33927;
	assign w33918 = w33929 & w33970;
	assign w33896 = w47755 ^ w44793;
	assign w33936 = w33896 ^ w33859;
	assign w33849 = w33896 ^ w33857;
	assign w33856 = w33886 ^ w33849;
	assign w33932 = w33853 ^ w33856;
	assign w33928 = w33849 ^ w33850;
	assign w33926 = w33936 & w33965;
	assign w33920 = w33928 & w33961;
	assign w33905 = w33920 ^ w44791;
	assign w33881 = w33920 ^ w33923;
	assign w33878 = ~w33881;
	assign w33877 = w33920 ^ w33921;
	assign w33871 = w33916 ^ w33905;
	assign w33868 = ~w33871;
	assign w33865 = w33921 ^ w33905;
	assign w33919 = w33932 & w33964;
	assign w33897 = w33915 ^ w33919;
	assign w33875 = ~w33897;
	assign w33874 = w33875 ^ w33913;
	assign w33870 = w33874 ^ w44792;
	assign w33873 = w33912 ^ w33870;
	assign w33917 = w33936 & w33967;
	assign w33911 = w33928 & w33976;
	assign w33910 = w33932 & w33973;
	assign w33876 = w33921 ^ w33910;
	assign w33872 = ~w33876;
	assign w33977 = w33872 ^ w33873;
	assign w48683 = ~w33977;
	assign w6495 = w45479 ^ w33977;
	assign w44790 = w33911 ^ w33912;
	assign w33893 = w33917 ^ w44790;
	assign w33894 = w33918 ^ w33893;
	assign w48685 = w33894 ^ w33865;
	assign w33898 = w33926 ^ w33894;
	assign w33867 = w33925 ^ w33898;
	assign w48681 = w33866 ^ w33867;
	assign w33903 = w33927 ^ w33898;
	assign w48682 = w44791 ^ w33903;
	assign w6674 = w48685 ^ w48689;
	assign w6455 = ~w6674;
	assign w6447 = ~w48681;
	assign w6457 = w48687 ^ w6447;
	assign w33978 = w33903 ^ w33877;
	assign w48684 = ~w33978;
	assign w6498 = w48688 ^ w48682;
	assign w6493 = w45480 ^ w33978;
	assign w33869 = w33893 ^ w33870;
	assign w48680 = w33868 ^ w33869;
	assign w6454 = ~w48680;
	assign w6453 = w48686 ^ w6454;
	assign w33880 = w33884 ^ w44790;
	assign w33883 = w44792 ^ w33880;
	assign w33980 = w33882 ^ w33883;
	assign w33879 = w33875 ^ w33880;
	assign w33979 = w33878 ^ w33879;
	assign w48679 = ~w33979;
	assign w6500 = w45481 ^ w33979;
	assign w45750 = ~w32369;
	assign w6550 = w6687 ^ w45750;
	assign w6684 = w45750 ^ w45566;
	assign w6580 = w6684 ^ w48673;
	assign w45751 = ~w32370;
	assign w6533 = w48670 ^ w45751;
	assign w45752 = ~w32371;
	assign w6702 = w45752 ^ w45568;
	assign w6547 = w6668 ^ w45752;
	assign w45753 = ~w32372;
	assign w6706 = w45753 ^ w45569;
	assign w6584 = w6706 ^ w6678;
	assign w45785 = ~w33980;
	assign w6451 = w45474 ^ w45785;
	assign w45804 = ~w38667;
	assign w48434 = w45804 ^ w6077;
	assign w6055 = w38668 ^ w45804;
	assign w6057 = w6056 ^ w6055;
	assign w48419 = ~w6057;
	assign w5999 = w45804 ^ w45488;
	assign w6065 = w5999 ^ w48504;
	assign w6041 = w5999 ^ w6011;
	assign w48411 = w45181 ^ w6041;
	assign w48426 = w6065 ^ w6064;
	assign w6052 = w5968 ^ w5999;
	assign w48418 = w45496 ^ w6052;
	assign w47654 = w48419 ^ w110;
	assign w34428 = w47660 ^ w47654;
	assign w47639 = w48434 ^ w125;
	assign w32010 = w47639 ^ w47637;
	assign w32085 = w32010 ^ w32100;
	assign w32093 = w32010 ^ w32016;
	assign w32096 = w47639 ^ w32016;
	assign w31972 = w32012 ^ w32010;
	assign w31971 = w32012 ^ w47639;
	assign w32095 = w47644 ^ w31971;
	assign w32081 = w47644 & w32095;
	assign w32076 = w32100 & w32085;
	assign w47655 = w48418 ^ w109;
	assign w34422 = w47655 ^ w47653;
	assign w34505 = w34422 ^ w34428;
	assign w34508 = w47655 ^ w34428;
	assign w47647 = w48426 ^ w117;
	assign w20754 = w47647 ^ w47645;
	assign w20829 = w20754 ^ w20844;
	assign w20837 = w20754 ^ w20760;
	assign w20840 = w47647 ^ w20760;
	assign w20716 = w20756 ^ w20754;
	assign w20715 = w20756 ^ w47647;
	assign w20839 = w47652 ^ w20715;
	assign w20825 = w47652 & w20839;
	assign w20820 = w20844 & w20829;
	assign w47662 = w48411 ^ w102;
	assign w20890 = w47664 ^ w47662;
	assign w20894 = w47668 ^ w47662;
	assign w20974 = w47663 ^ w20894;
	assign w20970 = w47667 ^ w20974;
	assign w20849 = w20890 ^ w47663;
	assign w20973 = w47668 ^ w20849;
	assign w20959 = w47668 & w20973;
	assign w20957 = w20974 & w20970;
	assign w45805 = ~w38669;
	assign w5979 = w45805 ^ w45182;
	assign w6070 = ~w5979;
	assign w6072 = w6070 ^ w5984;
	assign w48422 = w5939 ^ w5979;
	assign w47651 = w48422 ^ w113;
	assign w20753 = w47651 ^ w47649;
	assign w20755 = w47650 ^ w20753;
	assign w20831 = w47646 ^ w20755;
	assign w20828 = w47647 ^ w20755;
	assign w20830 = w20760 ^ w20755;
	assign w20836 = w47651 ^ w20840;
	assign w20834 = w20753 ^ w20842;
	assign w20833 = w47652 ^ w20834;
	assign w20770 = w47651 ^ w47650;
	assign w20835 = w20770 ^ w20837;
	assign w20838 = w20842 ^ w20770;
	assign w20832 = w20753 ^ w20716;
	assign w20843 = w47645 ^ w47651;
	assign w20827 = w20834 & w20838;
	assign w20759 = w20827 ^ w20756;
	assign w20826 = w20835 & w20833;
	assign w20777 = w20820 ^ w20826;
	assign w20824 = w20843 & w20828;
	assign w20758 = w20824 ^ w20754;
	assign w20823 = w20840 & w20836;
	assign w20822 = w20837 & w20830;
	assign w20821 = w20842 & w20831;
	assign w20757 = w20821 ^ w20755;
	assign w20763 = w20759 ^ w20757;
	assign w20768 = w47645 ^ w20763;
	assign w20818 = w20777 ^ w20768;
	assign w20729 = w20820 ^ w20821;
	assign w20776 = w20729 ^ w20730;
	assign w20775 = w20776 ^ w20758;
	assign w20817 = w20823 ^ w20775;
	assign w20819 = w20841 & w20832;
	assign w20814 = w20818 & w20817;
	assign w6048 = w5979 ^ w6016;
	assign w48415 = w48493 ^ w6048;
	assign w6225 = w6016 ^ w45805;
	assign w48407 = w6225 ^ w6224;
	assign w47666 = w48407 ^ w98;
	assign w20889 = w47666 ^ w20887;
	assign w20965 = w47662 ^ w20889;
	assign w20962 = w47663 ^ w20889;
	assign w20964 = w20894 ^ w20889;
	assign w20904 = w47667 ^ w47666;
	assign w20978 = w47666 ^ w47664;
	assign w20864 = w47665 ^ w47666;
	assign w47658 = w48415 ^ w106;
	assign w34509 = w47653 ^ w47658;
	assign w44238 = w20819 ^ w20825;
	assign w20731 = w20763 ^ w44238;
	assign w20774 = w47647 ^ w20731;
	assign w20809 = w20814 ^ w20774;
	assign w20769 = w44238 ^ w20754;
	assign w20815 = w20777 ^ w20769;
	assign w44239 = w20819 ^ w20822;
	assign w20772 = w20820 ^ w44239;
	assign w20728 = w20823 ^ w20772;
	assign w20810 = w47651 ^ w20728;
	assign w20808 = w20809 & w20810;
	assign w20806 = w20814 ^ w20808;
	assign w20727 = w20808 ^ w20772;
	assign w20726 = w20808 ^ w20825;
	assign w20721 = w20726 ^ w20822;
	assign w20732 = w20758 ^ w44239;
	assign w20816 = w20732 ^ w20757;
	assign w20807 = w20808 ^ w20816;
	assign w20813 = w20814 ^ w20816;
	assign w20812 = w20815 & w20813;
	assign w20811 = w20812 ^ w20774;
	assign w20723 = w20812 ^ w20824;
	assign w20719 = w20723 ^ w20759;
	assign w20722 = w47645 ^ w20719;
	assign w20799 = w20721 ^ w20722;
	assign w20720 = w20812 ^ w20768;
	assign w20718 = w47647 ^ w20719;
	assign w20805 = w20816 & w20806;
	assign w20803 = w20805 ^ w20813;
	assign w20802 = w20811 & w20803;
	assign w20767 = w20802 ^ w20777;
	assign w20801 = w20767 ^ w20769;
	assign w20725 = w20802 ^ w20826;
	assign w20798 = w20767 ^ w20720;
	assign w20793 = w20807 & w47652;
	assign w20792 = w20798 & w20828;
	assign w20791 = w20801 & w20840;
	assign w20790 = w20811 & w20830;
	assign w20734 = w20790 ^ w20791;
	assign w20789 = w20799 & w20831;
	assign w20784 = w20807 & w20839;
	assign w20783 = w20798 & w20843;
	assign w20750 = w20792 ^ w20783;
	assign w20782 = w20801 & w20836;
	assign w20752 = w20790 ^ w20782;
	assign w20781 = w20811 & w20837;
	assign w20780 = w20799 & w20842;
	assign w44241 = w20791 ^ w20792;
	assign w44243 = w20805 ^ w20823;
	assign w20797 = w44243 ^ w20775;
	assign w20795 = w20797 & w20834;
	assign w44242 = w20793 ^ w20795;
	assign w20786 = w20797 & w20838;
	assign w20764 = w47651 ^ w44243;
	assign w20804 = w20764 ^ w20727;
	assign w20717 = w20764 ^ w20725;
	assign w20724 = w20754 ^ w20717;
	assign w20800 = w20721 ^ w20724;
	assign w20796 = w20717 ^ w20718;
	assign w20794 = w20804 & w20833;
	assign w20788 = w20796 & w20829;
	assign w20773 = w20788 ^ w44241;
	assign w20749 = w20788 ^ w20791;
	assign w20746 = ~w20749;
	assign w20745 = w20788 ^ w20789;
	assign w20739 = w20784 ^ w20773;
	assign w20736 = ~w20739;
	assign w20733 = w20789 ^ w20773;
	assign w20787 = w20800 & w20832;
	assign w20765 = w20783 ^ w20787;
	assign w20743 = ~w20765;
	assign w20742 = w20743 ^ w20781;
	assign w20738 = w20742 ^ w44242;
	assign w20741 = w20780 ^ w20738;
	assign w20785 = w20804 & w20835;
	assign w20779 = w20796 & w20844;
	assign w20778 = w20800 & w20841;
	assign w20744 = w20789 ^ w20778;
	assign w20740 = ~w20744;
	assign w20845 = w20740 ^ w20741;
	assign w44240 = w20779 ^ w20780;
	assign w20761 = w20785 ^ w44240;
	assign w20737 = w20761 ^ w20738;
	assign w48649 = w20736 ^ w20737;
	assign w20762 = w20786 ^ w20761;
	assign w48652 = w20762 ^ w20733;
	assign w20766 = w20794 ^ w20762;
	assign w20735 = w20793 ^ w20766;
	assign w48650 = w20734 ^ w20735;
	assign w20771 = w20795 ^ w20766;
	assign w20846 = w20771 ^ w20745;
	assign w6468 = ~w48649;
	assign w6646 = w45657 ^ w6468;
	assign w6467 = w48650 ^ w6468;
	assign w48651 = w44241 ^ w20771;
	assign w20748 = w20752 ^ w44240;
	assign w20751 = w44242 ^ w20748;
	assign w20848 = w20750 ^ w20751;
	assign w20747 = w20743 ^ w20748;
	assign w20847 = w20746 ^ w20747;
	assign w48648 = ~w20847;
	assign w6461 = w20847 ^ w45650;
	assign w45467 = ~w20845;
	assign w45468 = ~w20846;
	assign w45469 = ~w20848;
	assign w6465 = w45657 ^ w45469;
	assign w45889 = ~w6029;
	assign w6207 = w45889 ^ w48492;
	assign w48396 = w6207 ^ w6206;
	assign w6184 = w45889 ^ w45486;
	assign w6186 = w6185 ^ w6184;
	assign w48382 = ~w6186;
	assign w47691 = w48382 ^ w73;
	assign w6411 = w47685 ^ w47691;
	assign w6338 = w47691 ^ w47690;
	assign w6188 = w45889 ^ w48475;
	assign w48384 = w6189 ^ w6188;
	assign w6190 = w45889 ^ w48476;
	assign w48385 = w6191 ^ w6190;
	assign w6403 = w6338 ^ w6405;
	assign w47688 = w48385 ^ w76;
	assign w6324 = w47688 ^ w47686;
	assign w6284 = w6324 ^ w6322;
	assign w6410 = w47688 ^ w47685;
	assign w6406 = w6410 ^ w6338;
	assign w6283 = w6324 ^ w47687;
	assign w6407 = w47692 ^ w6283;
	assign w6412 = w47690 ^ w47688;
	assign w6393 = w47692 & w6407;
	assign w47689 = w48384 ^ w75;
	assign w6321 = w47691 ^ w47689;
	assign w6400 = w6321 ^ w6284;
	assign w6402 = w6321 ^ w6410;
	assign w6395 = w6402 & w6406;
	assign w6327 = w6395 ^ w6324;
	assign w6401 = w47692 ^ w6402;
	assign w6394 = w6403 & w6401;
	assign w6387 = w6409 & w6400;
	assign w47677 = w48396 ^ w87;
	assign w25578 = w47679 ^ w47677;
	assign w25653 = w25578 ^ w25668;
	assign w25666 = w47680 ^ w47677;
	assign w25662 = w25666 ^ w25594;
	assign w25661 = w25578 ^ w25584;
	assign w25659 = w25594 ^ w25661;
	assign w25658 = w25577 ^ w25666;
	assign w25657 = w47684 ^ w25658;
	assign w25540 = w25580 ^ w25578;
	assign w25656 = w25577 ^ w25540;
	assign w25667 = w47677 ^ w47683;
	assign w25665 = w47677 ^ w47682;
	assign w25651 = w25658 & w25662;
	assign w25583 = w25651 ^ w25580;
	assign w25650 = w25659 & w25657;
	assign w25648 = w25667 & w25652;
	assign w25582 = w25648 ^ w25578;
	assign w25646 = w25661 & w25654;
	assign w25645 = w25666 & w25655;
	assign w25581 = w25645 ^ w25579;
	assign w25587 = w25583 ^ w25581;
	assign w25592 = w47677 ^ w25587;
	assign w25644 = w25668 & w25653;
	assign w25601 = w25644 ^ w25650;
	assign w25642 = w25601 ^ w25592;
	assign w25553 = w25644 ^ w25645;
	assign w25600 = w25553 ^ w25554;
	assign w25599 = w25600 ^ w25582;
	assign w25641 = w25647 ^ w25599;
	assign w25643 = w25665 & w25656;
	assign w25638 = w25642 & w25641;
	assign w6323 = w47690 ^ w6321;
	assign w6399 = w47686 ^ w6323;
	assign w6389 = w6410 & w6399;
	assign w6398 = w6328 ^ w6323;
	assign w6390 = w6405 & w6398;
	assign w6325 = w6389 ^ w6323;
	assign w6331 = w6327 ^ w6325;
	assign w6336 = w47685 ^ w6331;
	assign w6404 = w47691 ^ w6408;
	assign w6391 = w6408 & w6404;
	assign w6396 = w47687 ^ w6323;
	assign w6392 = w6411 & w6396;
	assign w6326 = w6392 ^ w6322;
	assign w43780 = w6387 ^ w6390;
	assign w6300 = w6326 ^ w43780;
	assign w6384 = w6300 ^ w6325;
	assign w43783 = w6387 ^ w6393;
	assign w6299 = w6331 ^ w43783;
	assign w6342 = w47687 ^ w6299;
	assign w6337 = w43783 ^ w6322;
	assign w44440 = w25643 ^ w25649;
	assign w25555 = w25587 ^ w44440;
	assign w25598 = w47679 ^ w25555;
	assign w25633 = w25638 ^ w25598;
	assign w25593 = w44440 ^ w25578;
	assign w25639 = w25601 ^ w25593;
	assign w44441 = w25643 ^ w25646;
	assign w25596 = w25644 ^ w44441;
	assign w25552 = w25647 ^ w25596;
	assign w25634 = w47683 ^ w25552;
	assign w25632 = w25633 & w25634;
	assign w25630 = w25638 ^ w25632;
	assign w25551 = w25632 ^ w25596;
	assign w25550 = w25632 ^ w25649;
	assign w25545 = w25550 ^ w25646;
	assign w25556 = w25582 ^ w44441;
	assign w25640 = w25556 ^ w25581;
	assign w25631 = w25632 ^ w25640;
	assign w25637 = w25638 ^ w25640;
	assign w25636 = w25639 & w25637;
	assign w25635 = w25636 ^ w25598;
	assign w25547 = w25636 ^ w25648;
	assign w25543 = w25547 ^ w25583;
	assign w25546 = w47677 ^ w25543;
	assign w25623 = w25545 ^ w25546;
	assign w25544 = w25636 ^ w25592;
	assign w25542 = w47679 ^ w25543;
	assign w25629 = w25640 & w25630;
	assign w25627 = w25629 ^ w25637;
	assign w25626 = w25635 & w25627;
	assign w25591 = w25626 ^ w25601;
	assign w25625 = w25591 ^ w25593;
	assign w25549 = w25626 ^ w25650;
	assign w25622 = w25591 ^ w25544;
	assign w25617 = w25631 & w47684;
	assign w25616 = w25622 & w25652;
	assign w25615 = w25625 & w25664;
	assign w25614 = w25635 & w25654;
	assign w25558 = w25614 ^ w25615;
	assign w25613 = w25623 & w25655;
	assign w25608 = w25631 & w25663;
	assign w25607 = w25622 & w25667;
	assign w25574 = w25616 ^ w25607;
	assign w25606 = w25625 & w25660;
	assign w25576 = w25614 ^ w25606;
	assign w25605 = w25635 & w25661;
	assign w25604 = w25623 & w25666;
	assign w44443 = w25615 ^ w25616;
	assign w44445 = w25629 ^ w25647;
	assign w25621 = w44445 ^ w25599;
	assign w25619 = w25621 & w25658;
	assign w44444 = w25617 ^ w25619;
	assign w25610 = w25621 & w25662;
	assign w25588 = w47683 ^ w44445;
	assign w25628 = w25588 ^ w25551;
	assign w25541 = w25588 ^ w25549;
	assign w25548 = w25578 ^ w25541;
	assign w25624 = w25545 ^ w25548;
	assign w25620 = w25541 ^ w25542;
	assign w25618 = w25628 & w25657;
	assign w25612 = w25620 & w25653;
	assign w25597 = w25612 ^ w44443;
	assign w25573 = w25612 ^ w25615;
	assign w25570 = ~w25573;
	assign w25569 = w25612 ^ w25613;
	assign w25563 = w25608 ^ w25597;
	assign w25560 = ~w25563;
	assign w25557 = w25613 ^ w25597;
	assign w25611 = w25624 & w25656;
	assign w25589 = w25607 ^ w25611;
	assign w25567 = ~w25589;
	assign w25566 = w25567 ^ w25605;
	assign w25562 = w25566 ^ w44444;
	assign w25565 = w25604 ^ w25562;
	assign w25609 = w25628 & w25659;
	assign w25603 = w25620 & w25668;
	assign w25602 = w25624 & w25665;
	assign w25568 = w25613 ^ w25602;
	assign w25564 = ~w25568;
	assign w25669 = w25564 ^ w25565;
	assign w44442 = w25603 ^ w25604;
	assign w25585 = w25609 ^ w44442;
	assign w25561 = w25585 ^ w25562;
	assign w48703 = w25560 ^ w25561;
	assign w25586 = w25610 ^ w25585;
	assign w48706 = w25586 ^ w25557;
	assign w25590 = w25618 ^ w25586;
	assign w25559 = w25617 ^ w25590;
	assign w48704 = w25558 ^ w25559;
	assign w25595 = w25619 ^ w25590;
	assign w25670 = w25595 ^ w25569;
	assign w48705 = w44443 ^ w25595;
	assign w6473 = w48705 ^ w48704;
	assign w25572 = w25576 ^ w44442;
	assign w25575 = w44444 ^ w25572;
	assign w25672 = w25574 ^ w25575;
	assign w25571 = w25567 ^ w25572;
	assign w25671 = w25570 ^ w25571;
	assign w6298 = w47689 ^ w47690;
	assign w6397 = w6322 ^ w6412;
	assign w6388 = w6412 & w6397;
	assign w6297 = w6388 ^ w6389;
	assign w6344 = w6297 ^ w6298;
	assign w6343 = w6344 ^ w6326;
	assign w6385 = w6391 ^ w6343;
	assign w6340 = w6388 ^ w43780;
	assign w6296 = w6391 ^ w6340;
	assign w6378 = w47691 ^ w6296;
	assign w6345 = w6388 ^ w6394;
	assign w6386 = w6345 ^ w6336;
	assign w6382 = w6386 & w6385;
	assign w6381 = w6382 ^ w6384;
	assign w6377 = w6382 ^ w6342;
	assign w6376 = w6377 & w6378;
	assign w6295 = w6376 ^ w6340;
	assign w6374 = w6382 ^ w6376;
	assign w6373 = w6384 & w6374;
	assign w6371 = w6373 ^ w6381;
	assign w6375 = w6376 ^ w6384;
	assign w6361 = w6375 & w47692;
	assign w6352 = w6375 & w6407;
	assign w43782 = w6373 ^ w6391;
	assign w6365 = w43782 ^ w6343;
	assign w6363 = w6365 & w6402;
	assign w6354 = w6365 & w6406;
	assign w6332 = w47691 ^ w43782;
	assign w6372 = w6332 ^ w6295;
	assign w6362 = w6372 & w6401;
	assign w6353 = w6372 & w6403;
	assign w43785 = w6361 ^ w6363;
	assign w6294 = w6376 ^ w6393;
	assign w6289 = w6294 ^ w6390;
	assign w6383 = w6345 ^ w6337;
	assign w6380 = w6383 & w6381;
	assign w6288 = w6380 ^ w6336;
	assign w6291 = w6380 ^ w6392;
	assign w6287 = w6291 ^ w6327;
	assign w6290 = w47685 ^ w6287;
	assign w6367 = w6289 ^ w6290;
	assign w6348 = w6367 & w6410;
	assign w6286 = w47687 ^ w6287;
	assign w6357 = w6367 & w6399;
	assign w6379 = w6380 ^ w6342;
	assign w6358 = w6379 & w6398;
	assign w6349 = w6379 & w6405;
	assign w6370 = w6379 & w6371;
	assign w6335 = w6370 ^ w6345;
	assign w6366 = w6335 ^ w6288;
	assign w6351 = w6366 & w6411;
	assign w6360 = w6366 & w6396;
	assign w6293 = w6370 ^ w6394;
	assign w6285 = w6332 ^ w6293;
	assign w6364 = w6285 ^ w6286;
	assign w6356 = w6364 & w6397;
	assign w6313 = w6356 ^ w6357;
	assign w6292 = w6322 ^ w6285;
	assign w6368 = w6289 ^ w6292;
	assign w6346 = w6368 & w6409;
	assign w6312 = w6357 ^ w6346;
	assign w6308 = ~w6312;
	assign w6318 = w6360 ^ w6351;
	assign w6355 = w6368 & w6400;
	assign w6333 = w6351 ^ w6355;
	assign w6311 = ~w6333;
	assign w6310 = w6311 ^ w6349;
	assign w6306 = w6310 ^ w43785;
	assign w6309 = w6348 ^ w6306;
	assign w6413 = w6308 ^ w6309;
	assign w6347 = w6364 & w6412;
	assign w48645 = ~w6413;
	assign w6369 = w6335 ^ w6337;
	assign w6359 = w6369 & w6408;
	assign w6350 = w6369 & w6404;
	assign w6320 = w6358 ^ w6350;
	assign w6317 = w6356 ^ w6359;
	assign w6314 = ~w6317;
	assign w6302 = w6358 ^ w6359;
	assign w6724 = w45655 ^ w48645;
	assign w6599 = w45467 ^ w6413;
	assign w43781 = w6347 ^ w6348;
	assign w6329 = w6353 ^ w43781;
	assign w6330 = w6354 ^ w6329;
	assign w6334 = w6362 ^ w6330;
	assign w6339 = w6363 ^ w6334;
	assign w6414 = w6339 ^ w6313;
	assign w48646 = ~w6414;
	assign w6722 = w45656 ^ w48646;
	assign w6597 = w45468 ^ w6414;
	assign w6305 = w6329 ^ w6306;
	assign w6316 = w6320 ^ w43781;
	assign w6319 = w43785 ^ w6316;
	assign w6315 = w6311 ^ w6316;
	assign w6415 = w6314 ^ w6315;
	assign w6416 = w6318 ^ w6319;
	assign w43784 = w6359 ^ w6360;
	assign w48644 = w43784 ^ w6339;
	assign w6601 = w48651 ^ w48644;
	assign w6727 = w48640 ^ w48644;
	assign w6341 = w6356 ^ w43784;
	assign w6307 = w6352 ^ w6341;
	assign w6304 = ~w6307;
	assign w6301 = w6357 ^ w6341;
	assign w48647 = w6330 ^ w6301;
	assign w6672 = w48641 ^ w48647;
	assign w6673 = w48647 ^ w48652;
	assign w48642 = w6304 ^ w6305;
	assign w6607 = ~w6673;
	assign w6711 = w48642 ^ w48649;
	assign w6594 = ~w6711;
	assign w6592 = w6594 ^ w48638;
	assign w6462 = w6672 ^ w48639;
	assign w6463 = w48638 ^ w48642;
	assign w6741 = w6462 ^ w6463;
	assign w6303 = w6361 ^ w6334;
	assign w48643 = w6302 ^ w6303;
	assign w6736 = w48639 ^ w48643;
	assign w6618 = ~w6736;
	assign w6605 = w6736 ^ w6594;
	assign w6459 = w48650 ^ w48643;
	assign w45191 = ~w6415;
	assign w6611 = w6607 ^ w45191;
	assign w6713 = w45191 ^ w48648;
	assign w45192 = ~w6416;
	assign w6712 = w45192 ^ w45469;
	assign w45562 = ~w25669;
	assign w45563 = ~w25670;
	assign w6621 = w45563 ^ w45562;
	assign w45564 = ~w25671;
	assign w45565 = ~w25672;
	assign w45900 = ~w6034;
	assign w6074 = w45900 ^ w48494;
	assign w6071 = w45900 ^ w45490;
	assign w6076 = w6075 ^ w6074;
	assign w48432 = ~w6076;
	assign w48430 = w6072 ^ w6071;
	assign w47643 = w48430 ^ w121;
	assign w32092 = w47643 ^ w32096;
	assign w32026 = w47643 ^ w47642;
	assign w32091 = w32026 ^ w32093;
	assign w32094 = w32098 ^ w32026;
	assign w32099 = w47637 ^ w47643;
	assign w32079 = w32096 & w32092;
	assign w6043 = w45900 ^ w45489;
	assign w48412 = w6043 ^ w6042;
	assign w47661 = w48412 ^ w103;
	assign w20888 = w47663 ^ w47661;
	assign w20963 = w20888 ^ w20978;
	assign w20976 = w47664 ^ w47661;
	assign w20972 = w20976 ^ w20904;
	assign w20971 = w20888 ^ w20894;
	assign w20969 = w20904 ^ w20971;
	assign w20968 = w20887 ^ w20976;
	assign w20967 = w47668 ^ w20968;
	assign w20850 = w20890 ^ w20888;
	assign w20966 = w20887 ^ w20850;
	assign w20977 = w47661 ^ w47667;
	assign w20975 = w47661 ^ w47666;
	assign w20961 = w20968 & w20972;
	assign w20893 = w20961 ^ w20890;
	assign w20960 = w20969 & w20967;
	assign w20958 = w20977 & w20962;
	assign w20892 = w20958 ^ w20888;
	assign w20956 = w20971 & w20964;
	assign w20955 = w20976 & w20965;
	assign w20891 = w20955 ^ w20889;
	assign w20897 = w20893 ^ w20891;
	assign w20902 = w47661 ^ w20897;
	assign w20954 = w20978 & w20963;
	assign w20911 = w20954 ^ w20960;
	assign w20952 = w20911 ^ w20902;
	assign w20863 = w20954 ^ w20955;
	assign w20910 = w20863 ^ w20864;
	assign w20909 = w20910 ^ w20892;
	assign w20951 = w20957 ^ w20909;
	assign w20953 = w20975 & w20966;
	assign w20948 = w20952 & w20951;
	assign w44244 = w20953 ^ w20959;
	assign w20903 = w44244 ^ w20888;
	assign w20949 = w20911 ^ w20903;
	assign w20865 = w20897 ^ w44244;
	assign w20908 = w47663 ^ w20865;
	assign w20943 = w20948 ^ w20908;
	assign w44245 = w20953 ^ w20956;
	assign w20906 = w20954 ^ w44245;
	assign w20862 = w20957 ^ w20906;
	assign w20944 = w47667 ^ w20862;
	assign w20942 = w20943 & w20944;
	assign w20861 = w20942 ^ w20906;
	assign w20860 = w20942 ^ w20959;
	assign w20855 = w20860 ^ w20956;
	assign w20940 = w20948 ^ w20942;
	assign w20866 = w20892 ^ w44245;
	assign w20950 = w20866 ^ w20891;
	assign w20941 = w20942 ^ w20950;
	assign w20947 = w20948 ^ w20950;
	assign w20946 = w20949 & w20947;
	assign w20945 = w20946 ^ w20908;
	assign w20857 = w20946 ^ w20958;
	assign w20853 = w20857 ^ w20893;
	assign w20856 = w47661 ^ w20853;
	assign w20933 = w20855 ^ w20856;
	assign w20854 = w20946 ^ w20902;
	assign w20852 = w47663 ^ w20853;
	assign w20939 = w20950 & w20940;
	assign w20937 = w20939 ^ w20947;
	assign w20936 = w20945 & w20937;
	assign w20901 = w20936 ^ w20911;
	assign w20935 = w20901 ^ w20903;
	assign w20859 = w20936 ^ w20960;
	assign w20932 = w20901 ^ w20854;
	assign w20927 = w20941 & w47668;
	assign w20926 = w20932 & w20962;
	assign w20925 = w20935 & w20974;
	assign w20924 = w20945 & w20964;
	assign w20868 = w20924 ^ w20925;
	assign w20923 = w20933 & w20965;
	assign w20918 = w20941 & w20973;
	assign w20917 = w20932 & w20977;
	assign w20884 = w20926 ^ w20917;
	assign w20916 = w20935 & w20970;
	assign w20886 = w20924 ^ w20916;
	assign w20915 = w20945 & w20971;
	assign w20914 = w20933 & w20976;
	assign w44246 = w20925 ^ w20926;
	assign w44248 = w20939 ^ w20957;
	assign w20898 = w47667 ^ w44248;
	assign w20938 = w20898 ^ w20861;
	assign w20919 = w20938 & w20969;
	assign w20928 = w20938 & w20967;
	assign w20851 = w20898 ^ w20859;
	assign w20858 = w20888 ^ w20851;
	assign w20934 = w20855 ^ w20858;
	assign w20921 = w20934 & w20966;
	assign w20899 = w20917 ^ w20921;
	assign w20877 = ~w20899;
	assign w20876 = w20877 ^ w20915;
	assign w20930 = w20851 ^ w20852;
	assign w20913 = w20930 & w20978;
	assign w20912 = w20934 & w20975;
	assign w20878 = w20923 ^ w20912;
	assign w20874 = ~w20878;
	assign w43557 = w20913 ^ w20914;
	assign w20895 = w20919 ^ w43557;
	assign w20882 = w20886 ^ w43557;
	assign w20881 = w20877 ^ w20882;
	assign w20922 = w20930 & w20963;
	assign w20879 = w20922 ^ w20923;
	assign w20907 = w20922 ^ w44246;
	assign w20873 = w20918 ^ w20907;
	assign w20870 = ~w20873;
	assign w20867 = w20923 ^ w20907;
	assign w20883 = w20922 ^ w20925;
	assign w20880 = ~w20883;
	assign w20981 = w20880 ^ w20881;
	assign w20931 = w44248 ^ w20909;
	assign w20929 = w20931 & w20968;
	assign w20920 = w20931 & w20972;
	assign w20896 = w20920 ^ w20895;
	assign w20900 = w20928 ^ w20896;
	assign w20905 = w20929 ^ w20900;
	assign w48677 = w44246 ^ w20905;
	assign w20980 = w20905 ^ w20879;
	assign w20869 = w20927 ^ w20900;
	assign w48676 = w20868 ^ w20869;
	assign w48678 = w20896 ^ w20867;
	assign w6670 = w48678 ^ w48685;
	assign w6710 = w48677 ^ w48682;
	assign w6718 = w48676 ^ w48681;
	assign w6526 = w33977 ^ w48677;
	assign w6482 = ~w6710;
	assign w6485 = ~w6718;
	assign w6449 = w48682 ^ w48676;
	assign w44247 = w20927 ^ w20929;
	assign w20885 = w44247 ^ w20882;
	assign w20982 = w20884 ^ w20885;
	assign w20872 = w20876 ^ w44247;
	assign w20875 = w20914 ^ w20872;
	assign w20979 = w20874 ^ w20875;
	assign w20871 = w20895 ^ w20872;
	assign w48675 = w20870 ^ w20871;
	assign w6725 = w48675 ^ w48680;
	assign w6501 = ~w6725;
	assign w6446 = w6447 ^ w48675;
	assign w47641 = w48432 ^ w123;
	assign w32009 = w47643 ^ w47641;
	assign w32011 = w47642 ^ w32009;
	assign w32087 = w47638 ^ w32011;
	assign w32084 = w47639 ^ w32011;
	assign w32086 = w32016 ^ w32011;
	assign w32090 = w32009 ^ w32098;
	assign w32089 = w47644 ^ w32090;
	assign w31986 = w47641 ^ w47642;
	assign w32088 = w32009 ^ w31972;
	assign w32083 = w32090 & w32094;
	assign w32015 = w32083 ^ w32012;
	assign w32082 = w32091 & w32089;
	assign w32033 = w32076 ^ w32082;
	assign w32080 = w32099 & w32084;
	assign w32014 = w32080 ^ w32010;
	assign w32078 = w32093 & w32086;
	assign w32077 = w32098 & w32087;
	assign w32013 = w32077 ^ w32011;
	assign w32019 = w32015 ^ w32013;
	assign w32024 = w47637 ^ w32019;
	assign w32074 = w32033 ^ w32024;
	assign w31985 = w32076 ^ w32077;
	assign w32032 = w31985 ^ w31986;
	assign w32031 = w32032 ^ w32014;
	assign w32073 = w32079 ^ w32031;
	assign w32075 = w32097 & w32088;
	assign w32070 = w32074 & w32073;
	assign w44711 = w32075 ^ w32078;
	assign w31988 = w32014 ^ w44711;
	assign w32072 = w31988 ^ w32013;
	assign w32069 = w32070 ^ w32072;
	assign w32028 = w32076 ^ w44711;
	assign w31984 = w32079 ^ w32028;
	assign w32066 = w47643 ^ w31984;
	assign w44714 = w32075 ^ w32081;
	assign w31987 = w32019 ^ w44714;
	assign w32030 = w47639 ^ w31987;
	assign w32065 = w32070 ^ w32030;
	assign w32064 = w32065 & w32066;
	assign w32062 = w32070 ^ w32064;
	assign w31983 = w32064 ^ w32028;
	assign w31982 = w32064 ^ w32081;
	assign w31977 = w31982 ^ w32078;
	assign w32061 = w32072 & w32062;
	assign w32059 = w32061 ^ w32069;
	assign w44713 = w32061 ^ w32079;
	assign w32053 = w44713 ^ w32031;
	assign w32042 = w32053 & w32094;
	assign w32051 = w32053 & w32090;
	assign w32020 = w47643 ^ w44713;
	assign w32060 = w32020 ^ w31983;
	assign w32050 = w32060 & w32089;
	assign w32041 = w32060 & w32091;
	assign w32063 = w32064 ^ w32072;
	assign w32049 = w32063 & w47644;
	assign w32040 = w32063 & w32095;
	assign w32025 = w44714 ^ w32010;
	assign w32071 = w32033 ^ w32025;
	assign w32068 = w32071 & w32069;
	assign w32067 = w32068 ^ w32030;
	assign w31979 = w32068 ^ w32080;
	assign w31975 = w31979 ^ w32015;
	assign w31978 = w47637 ^ w31975;
	assign w32055 = w31977 ^ w31978;
	assign w31976 = w32068 ^ w32024;
	assign w31974 = w47639 ^ w31975;
	assign w32058 = w32067 & w32059;
	assign w32023 = w32058 ^ w32033;
	assign w32057 = w32023 ^ w32025;
	assign w31981 = w32058 ^ w32082;
	assign w31973 = w32020 ^ w31981;
	assign w31980 = w32010 ^ w31973;
	assign w32056 = w31977 ^ w31980;
	assign w32054 = w32023 ^ w31976;
	assign w32052 = w31973 ^ w31974;
	assign w32048 = w32054 & w32084;
	assign w32047 = w32057 & w32096;
	assign w32046 = w32067 & w32086;
	assign w31990 = w32046 ^ w32047;
	assign w32045 = w32055 & w32087;
	assign w32044 = w32052 & w32085;
	assign w32005 = w32044 ^ w32047;
	assign w32002 = ~w32005;
	assign w32001 = w32044 ^ w32045;
	assign w32043 = w32056 & w32088;
	assign w32039 = w32054 & w32099;
	assign w32021 = w32039 ^ w32043;
	assign w32006 = w32048 ^ w32039;
	assign w31999 = ~w32021;
	assign w32038 = w32057 & w32092;
	assign w32008 = w32046 ^ w32038;
	assign w32037 = w32067 & w32093;
	assign w31998 = w31999 ^ w32037;
	assign w32036 = w32055 & w32098;
	assign w32035 = w32052 & w32100;
	assign w32034 = w32056 & w32097;
	assign w32000 = w32045 ^ w32034;
	assign w31996 = ~w32000;
	assign w44712 = w32035 ^ w32036;
	assign w32017 = w32041 ^ w44712;
	assign w32018 = w32042 ^ w32017;
	assign w32022 = w32050 ^ w32018;
	assign w31991 = w32049 ^ w32022;
	assign w48708 = w31990 ^ w31991;
	assign w32027 = w32051 ^ w32022;
	assign w32102 = w32027 ^ w32001;
	assign w32004 = w32008 ^ w44712;
	assign w32003 = w31999 ^ w32004;
	assign w32103 = w32002 ^ w32003;
	assign w44715 = w32047 ^ w32048;
	assign w48709 = w44715 ^ w32027;
	assign w6682 = w48705 ^ w48709;
	assign w32029 = w32044 ^ w44715;
	assign w31995 = w32040 ^ w32029;
	assign w31992 = ~w31995;
	assign w31989 = w32045 ^ w32029;
	assign w48710 = w32018 ^ w31989;
	assign w6665 = w48706 ^ w48710;
	assign w6472 = w6665 ^ w48708;
	assign w6737 = w6472 ^ w6473;
	assign w44716 = w32049 ^ w32051;
	assign w32007 = w44716 ^ w32004;
	assign w32104 = w32006 ^ w32007;
	assign w31994 = w31998 ^ w44716;
	assign w31997 = w32036 ^ w31994;
	assign w32101 = w31996 ^ w31997;
	assign w31993 = w32017 ^ w31994;
	assign w48707 = w31992 ^ w31993;
	assign w6683 = w48703 ^ w48707;
	assign w6434 = w48708 ^ w48707;
	assign w45466 = ~w20982;
	assign w6733 = w45466 ^ w45785;
	assign w6502 = w6733 ^ w6674;
	assign w6443 = w33979 ^ w45466;
	assign w45471 = ~w20979;
	assign w6703 = w45471 ^ w48683;
	assign w6521 = w33978 ^ w45471;
	assign w45472 = ~w20980;
	assign w6696 = w45472 ^ w48684;
	assign w6518 = w48685 ^ w45472;
	assign w45473 = ~w20981;
	assign w6732 = w45473 ^ w48679;
	assign w6529 = w6454 ^ w45473;
	assign w45742 = ~w32101;
	assign w45743 = ~w32102;
	assign w6688 = w45563 ^ w45743;
	assign w45744 = ~w32103;
	assign w6695 = w45564 ^ w45744;
	assign w45745 = ~w32104;
	assign w6715 = w45565 ^ w45745;
	assign w45888 = ~w6670;
	assign w6511 = w45888 ^ w48676;
	assign w6515 = w45888 ^ w45473;
	assign w6509 = w45888 ^ w48677;
	assign w45901 = ~w6028;
	assign w6109 = w45901 ^ w48450;
	assign w48337 = w6110 ^ w6109;
	assign w6196 = w45901 ^ w45505;
	assign w48316 = w6196 ^ w6195;
	assign w6233 = w45901 ^ w48452;
	assign w5960 = w6233 ^ w6232;
	assign w48336 = w5960 ^ w5963;
	assign w47736 = w48337 ^ w28;
	assign w21292 = w47736 ^ w47734;
	assign w21378 = w47736 ^ w47733;
	assign w21374 = w21378 ^ w21306;
	assign w21380 = w47738 ^ w47736;
	assign w21365 = w21290 ^ w21380;
	assign w21252 = w21292 ^ w21290;
	assign w21251 = w21292 ^ w47735;
	assign w21375 = w47740 ^ w21251;
	assign w21361 = w47740 & w21375;
	assign w21356 = w21380 & w21365;
	assign w47737 = w48336 ^ w27;
	assign w21289 = w47739 ^ w47737;
	assign w21291 = w47738 ^ w21289;
	assign w21367 = w47734 ^ w21291;
	assign w21364 = w47735 ^ w21291;
	assign w21366 = w21296 ^ w21291;
	assign w21370 = w21289 ^ w21378;
	assign w21369 = w47740 ^ w21370;
	assign w21266 = w47737 ^ w47738;
	assign w21368 = w21289 ^ w21252;
	assign w21363 = w21370 & w21374;
	assign w21295 = w21363 ^ w21292;
	assign w21362 = w21371 & w21369;
	assign w21313 = w21356 ^ w21362;
	assign w21360 = w21379 & w21364;
	assign w21294 = w21360 ^ w21290;
	assign w21358 = w21373 & w21366;
	assign w21357 = w21378 & w21367;
	assign w21293 = w21357 ^ w21291;
	assign w21299 = w21295 ^ w21293;
	assign w21304 = w47733 ^ w21299;
	assign w21354 = w21313 ^ w21304;
	assign w21265 = w21356 ^ w21357;
	assign w21312 = w21265 ^ w21266;
	assign w21311 = w21312 ^ w21294;
	assign w21353 = w21359 ^ w21311;
	assign w21355 = w21377 & w21368;
	assign w21350 = w21354 & w21353;
	assign w47757 = w48316 ^ w7;
	assign w32412 = w47759 ^ w47757;
	assign w32487 = w32412 ^ w32502;
	assign w32500 = w47760 ^ w47757;
	assign w32496 = w32500 ^ w32428;
	assign w32495 = w32412 ^ w32418;
	assign w32493 = w32428 ^ w32495;
	assign w32492 = w32411 ^ w32500;
	assign w32491 = w47764 ^ w32492;
	assign w32374 = w32414 ^ w32412;
	assign w32490 = w32411 ^ w32374;
	assign w32501 = w47757 ^ w47763;
	assign w32499 = w47757 ^ w47762;
	assign w32485 = w32492 & w32496;
	assign w32417 = w32485 ^ w32414;
	assign w32484 = w32493 & w32491;
	assign w32482 = w32501 & w32486;
	assign w32416 = w32482 ^ w32412;
	assign w32480 = w32495 & w32488;
	assign w32479 = w32500 & w32489;
	assign w32415 = w32479 ^ w32413;
	assign w32421 = w32417 ^ w32415;
	assign w32426 = w47757 ^ w32421;
	assign w32478 = w32502 & w32487;
	assign w32435 = w32478 ^ w32484;
	assign w32476 = w32435 ^ w32426;
	assign w32387 = w32478 ^ w32479;
	assign w32434 = w32387 ^ w32388;
	assign w32433 = w32434 ^ w32416;
	assign w32475 = w32481 ^ w32433;
	assign w32477 = w32499 & w32490;
	assign w32472 = w32476 & w32475;
	assign w44261 = w21355 ^ w21361;
	assign w21305 = w44261 ^ w21290;
	assign w21351 = w21313 ^ w21305;
	assign w21267 = w21299 ^ w44261;
	assign w21310 = w47735 ^ w21267;
	assign w21345 = w21350 ^ w21310;
	assign w44262 = w21355 ^ w21358;
	assign w21308 = w21356 ^ w44262;
	assign w21264 = w21359 ^ w21308;
	assign w21346 = w47739 ^ w21264;
	assign w21344 = w21345 & w21346;
	assign w21342 = w21350 ^ w21344;
	assign w21263 = w21344 ^ w21308;
	assign w21262 = w21344 ^ w21361;
	assign w21257 = w21262 ^ w21358;
	assign w21268 = w21294 ^ w44262;
	assign w21352 = w21268 ^ w21293;
	assign w21343 = w21344 ^ w21352;
	assign w21349 = w21350 ^ w21352;
	assign w21348 = w21351 & w21349;
	assign w21347 = w21348 ^ w21310;
	assign w21259 = w21348 ^ w21360;
	assign w21255 = w21259 ^ w21295;
	assign w21258 = w47733 ^ w21255;
	assign w21335 = w21257 ^ w21258;
	assign w21256 = w21348 ^ w21304;
	assign w21254 = w47735 ^ w21255;
	assign w21341 = w21352 & w21342;
	assign w21339 = w21341 ^ w21349;
	assign w21338 = w21347 & w21339;
	assign w21303 = w21338 ^ w21313;
	assign w21337 = w21303 ^ w21305;
	assign w21261 = w21338 ^ w21362;
	assign w21334 = w21303 ^ w21256;
	assign w21329 = w21343 & w47740;
	assign w21328 = w21334 & w21364;
	assign w21327 = w21337 & w21376;
	assign w21326 = w21347 & w21366;
	assign w21270 = w21326 ^ w21327;
	assign w21325 = w21335 & w21367;
	assign w21320 = w21343 & w21375;
	assign w21319 = w21334 & w21379;
	assign w21286 = w21328 ^ w21319;
	assign w21318 = w21337 & w21372;
	assign w21288 = w21326 ^ w21318;
	assign w21317 = w21347 & w21373;
	assign w21316 = w21335 & w21378;
	assign w44263 = w21327 ^ w21328;
	assign w44265 = w21341 ^ w21359;
	assign w21300 = w47739 ^ w44265;
	assign w21253 = w21300 ^ w21261;
	assign w21260 = w21290 ^ w21253;
	assign w21336 = w21257 ^ w21260;
	assign w21323 = w21336 & w21368;
	assign w21301 = w21319 ^ w21323;
	assign w21279 = ~w21301;
	assign w21332 = w21253 ^ w21254;
	assign w21324 = w21332 & w21365;
	assign w21285 = w21324 ^ w21327;
	assign w21282 = ~w21285;
	assign w21281 = w21324 ^ w21325;
	assign w21278 = w21279 ^ w21317;
	assign w21315 = w21332 & w21380;
	assign w21314 = w21336 & w21377;
	assign w21280 = w21325 ^ w21314;
	assign w21276 = ~w21280;
	assign w43558 = w21315 ^ w21316;
	assign w21284 = w21288 ^ w43558;
	assign w21283 = w21279 ^ w21284;
	assign w21383 = w21282 ^ w21283;
	assign w21309 = w21324 ^ w44263;
	assign w21275 = w21320 ^ w21309;
	assign w21272 = ~w21275;
	assign w21269 = w21325 ^ w21309;
	assign w21340 = w21300 ^ w21263;
	assign w21321 = w21340 & w21371;
	assign w21297 = w21321 ^ w43558;
	assign w21330 = w21340 & w21369;
	assign w21333 = w44265 ^ w21311;
	assign w21331 = w21333 & w21370;
	assign w21322 = w21333 & w21374;
	assign w21298 = w21322 ^ w21297;
	assign w21302 = w21330 ^ w21298;
	assign w21307 = w21331 ^ w21302;
	assign w48655 = w44263 ^ w21307;
	assign w21382 = w21307 ^ w21281;
	assign w21271 = w21329 ^ w21302;
	assign w48654 = w21270 ^ w21271;
	assign w48657 = w21298 ^ w21269;
	assign w48656 = ~w21382;
	assign w6541 = w48655 ^ w6413;
	assign w6671 = w48652 ^ w48657;
	assign w6723 = w48651 ^ w48655;
	assign w6726 = w48650 ^ w48654;
	assign w48521 = w6741 ^ w6726;
	assign w47625 = w48521 ^ w1989;
	assign w6613 = w6722 ^ w6671;
	assign w6598 = w6722 ^ w21382;
	assign w48532 = w6598 ^ w6599;
	assign w47614 = w48532 ^ w2000;
	assign w6616 = w6618 ^ w6723;
	assign w6606 = w6607 ^ w48654;
	assign w6716 = w45468 ^ w48656;
	assign w6614 = w6724 ^ w6716;
	assign w6585 = w6716 ^ w6672;
	assign w48524 = w45656 ^ w6614;
	assign w47622 = w48524 ^ w1992;
	assign w48525 = w48641 ^ w6613;
	assign w47621 = w48525 ^ w1993;
	assign w48529 = w6605 ^ w6606;
	assign w47617 = w48529 ^ w1997;
	assign w6595 = w6712 ^ w6671;
	assign w6458 = w6673 ^ w48655;
	assign w6743 = w6458 ^ w6459;
	assign w48530 = w6743 ^ w6727;
	assign w47616 = w48530 ^ w1998;
	assign w20622 = w47616 ^ w47614;
	assign w6591 = w6727 ^ w6726;
	assign w6589 = ~w6591;
	assign w6523 = w6716 ^ w45655;
	assign w6504 = w21382 ^ w48647;
	assign w48541 = w48652 ^ w6585;
	assign w47605 = w48541 ^ w2009;
	assign w6679 = w48641 ^ w48657;
	assign w6664 = w6712 ^ w6679;
	assign w6575 = ~w6679;
	assign w6574 = w6575 ^ w48643;
	assign w48534 = w45650 ^ w6595;
	assign w47612 = w48534 ^ w2002;
	assign w6588 = w6724 ^ w6723;
	assign w6421 = w6679 ^ w48639;
	assign w6422 = w48654 ^ w48644;
	assign w6758 = w6421 ^ w6422;
	assign w48514 = w6758 ^ w6723;
	assign w47632 = w48514 ^ w1982;
	assign w44264 = w21329 ^ w21331;
	assign w21287 = w44264 ^ w21284;
	assign w21384 = w21286 ^ w21287;
	assign w21274 = w21278 ^ w44264;
	assign w21277 = w21316 ^ w21274;
	assign w21381 = w21276 ^ w21277;
	assign w21273 = w21297 ^ w21274;
	assign w48653 = w21272 ^ w21273;
	assign w6714 = w48638 ^ w48653;
	assign w6576 = ~w6714;
	assign w6573 = w6726 ^ w6576;
	assign w6608 = w6714 ^ w6713;
	assign w48528 = w48642 ^ w6608;
	assign w47618 = w48528 ^ w1996;
	assign w20710 = w47618 ^ w47616;
	assign w20596 = w47617 ^ w47618;
	assign w6645 = w6576 ^ w45191;
	assign w48520 = w6645 ^ w6646;
	assign w47626 = w48520 ^ w1988;
	assign w13896 = w47625 ^ w47626;
	assign w14007 = w47621 ^ w47626;
	assign w48513 = w6573 ^ w6574;
	assign w47633 = w48513 ^ w1981;
	assign w44727 = w32477 ^ w32480;
	assign w32390 = w32416 ^ w44727;
	assign w32474 = w32390 ^ w32415;
	assign w32471 = w32472 ^ w32474;
	assign w32430 = w32478 ^ w44727;
	assign w32386 = w32481 ^ w32430;
	assign w32468 = w47763 ^ w32386;
	assign w44730 = w32477 ^ w32483;
	assign w32389 = w32421 ^ w44730;
	assign w32432 = w47759 ^ w32389;
	assign w32467 = w32472 ^ w32432;
	assign w32466 = w32467 & w32468;
	assign w32464 = w32472 ^ w32466;
	assign w32385 = w32466 ^ w32430;
	assign w32384 = w32466 ^ w32483;
	assign w32379 = w32384 ^ w32480;
	assign w32463 = w32474 & w32464;
	assign w32461 = w32463 ^ w32471;
	assign w44729 = w32463 ^ w32481;
	assign w32455 = w44729 ^ w32433;
	assign w32444 = w32455 & w32496;
	assign w32453 = w32455 & w32492;
	assign w32422 = w47763 ^ w44729;
	assign w32462 = w32422 ^ w32385;
	assign w32452 = w32462 & w32491;
	assign w32443 = w32462 & w32493;
	assign w32465 = w32466 ^ w32474;
	assign w32451 = w32465 & w47764;
	assign w32442 = w32465 & w32497;
	assign w32427 = w44730 ^ w32412;
	assign w32473 = w32435 ^ w32427;
	assign w32470 = w32473 & w32471;
	assign w32469 = w32470 ^ w32432;
	assign w32381 = w32470 ^ w32482;
	assign w32377 = w32381 ^ w32417;
	assign w32380 = w47757 ^ w32377;
	assign w32457 = w32379 ^ w32380;
	assign w32378 = w32470 ^ w32426;
	assign w32376 = w47759 ^ w32377;
	assign w32460 = w32469 & w32461;
	assign w32425 = w32460 ^ w32435;
	assign w32459 = w32425 ^ w32427;
	assign w32383 = w32460 ^ w32484;
	assign w32375 = w32422 ^ w32383;
	assign w32382 = w32412 ^ w32375;
	assign w32458 = w32379 ^ w32382;
	assign w32456 = w32425 ^ w32378;
	assign w32454 = w32375 ^ w32376;
	assign w32450 = w32456 & w32486;
	assign w32449 = w32459 & w32498;
	assign w32448 = w32469 & w32488;
	assign w32392 = w32448 ^ w32449;
	assign w32447 = w32457 & w32489;
	assign w32446 = w32454 & w32487;
	assign w32407 = w32446 ^ w32449;
	assign w32404 = ~w32407;
	assign w32403 = w32446 ^ w32447;
	assign w32445 = w32458 & w32490;
	assign w32441 = w32456 & w32501;
	assign w32423 = w32441 ^ w32445;
	assign w32408 = w32450 ^ w32441;
	assign w32401 = ~w32423;
	assign w32440 = w32459 & w32494;
	assign w32410 = w32448 ^ w32440;
	assign w32439 = w32469 & w32495;
	assign w32400 = w32401 ^ w32439;
	assign w32438 = w32457 & w32500;
	assign w32437 = w32454 & w32502;
	assign w32436 = w32458 & w32499;
	assign w32402 = w32447 ^ w32436;
	assign w32398 = ~w32402;
	assign w44728 = w32437 ^ w32438;
	assign w32419 = w32443 ^ w44728;
	assign w32420 = w32444 ^ w32419;
	assign w32424 = w32452 ^ w32420;
	assign w32393 = w32451 ^ w32424;
	assign w48695 = w32392 ^ w32393;
	assign w6691 = w48695 ^ w48708;
	assign w6662 = w6691 ^ w6682;
	assign w32429 = w32453 ^ w32424;
	assign w32504 = w32429 ^ w32403;
	assign w48697 = ~w32504;
	assign w32406 = w32410 ^ w44728;
	assign w32405 = w32401 ^ w32406;
	assign w32505 = w32404 ^ w32405;
	assign w44731 = w32449 ^ w32450;
	assign w48696 = w44731 ^ w32429;
	assign w6471 = ~w48696;
	assign w6660 = w48709 ^ w6471;
	assign w32431 = w32446 ^ w44731;
	assign w32397 = w32442 ^ w32431;
	assign w32394 = ~w32397;
	assign w32391 = w32447 ^ w32431;
	assign w48698 = w32420 ^ w32391;
	assign w6677 = w48698 ^ w48710;
	assign w6476 = w6715 ^ w6677;
	assign w44732 = w32451 ^ w32453;
	assign w32409 = w44732 ^ w32406;
	assign w32506 = w32408 ^ w32409;
	assign w32396 = w32400 ^ w44732;
	assign w32399 = w32438 ^ w32396;
	assign w32503 = w32398 ^ w32399;
	assign w32395 = w32419 ^ w32396;
	assign w48694 = w32394 ^ w32395;
	assign w6433 = w6677 ^ w48694;
	assign w6753 = w6433 ^ w6434;
	assign w48539 = w45467 ^ w6588;
	assign w47607 = w48539 ^ w2007;
	assign w28660 = w47607 ^ w47605;
	assign w45478 = ~w21384;
	assign w6735 = w45650 ^ w45478;
	assign w6603 = w6735 ^ w6713;
	assign w6612 = w6735 ^ w6673;
	assign w48510 = w45478 ^ w6664;
	assign w47636 = w48510 ^ w1978;
	assign w48526 = w45192 ^ w6612;
	assign w47620 = w48526 ^ w1994;
	assign w20626 = w47620 ^ w47614;
	assign w6464 = w6671 ^ w45478;
	assign w6740 = w6464 ^ w6465;
	assign w6487 = w6735 ^ w6672;
	assign w48518 = w45469 ^ w6487;
	assign w47628 = w48518 ^ w1986;
	assign w13926 = w47628 ^ w47622;
	assign w48535 = w6740 ^ w6713;
	assign w47611 = w48535 ^ w2003;
	assign w28749 = w47605 ^ w47611;
	assign w45484 = ~w21381;
	assign w6600 = w6724 ^ w45484;
	assign w6524 = w45484 ^ w6414;
	assign w6522 = w6523 ^ w6524;
	assign w48516 = ~w6522;
	assign w47630 = w48516 ^ w1984;
	assign w25446 = w47632 ^ w47630;
	assign w25450 = w47636 ^ w47630;
	assign w48531 = w6600 ^ w6601;
	assign w47615 = w48531 ^ w1999;
	assign w20706 = w47615 ^ w20626;
	assign w20581 = w20622 ^ w47615;
	assign w20705 = w47620 ^ w20581;
	assign w20691 = w47620 & w20705;
	assign w6719 = w45467 ^ w45484;
	assign w6615 = w6727 ^ w6719;
	assign w48523 = w45655 ^ w6615;
	assign w47623 = w48523 ^ w1991;
	assign w13920 = w47623 ^ w47621;
	assign w14003 = w13920 ^ w13926;
	assign w14006 = w47623 ^ w13926;
	assign w6586 = w6722 ^ w6719;
	assign w48540 = w45468 ^ w6586;
	assign w47606 = w48540 ^ w2008;
	assign w28666 = w47612 ^ w47606;
	assign w28743 = w28660 ^ w28666;
	assign w28746 = w47607 ^ w28666;
	assign w28742 = w47611 ^ w28746;
	assign w28729 = w28746 & w28742;
	assign w6542 = w6719 ^ w48640;
	assign w6540 = ~w6542;
	assign w48515 = w6540 ^ w6541;
	assign w47631 = w48515 ^ w1983;
	assign w25530 = w47631 ^ w25450;
	assign w25405 = w25446 ^ w47631;
	assign w25529 = w47636 ^ w25405;
	assign w25515 = w47636 & w25529;
	assign w45485 = ~w21383;
	assign w6734 = w45657 ^ w45485;
	assign w6587 = w6734 ^ w6711;
	assign w48512 = w48653 ^ w6587;
	assign w47634 = w48512 ^ w1980;
	assign w25534 = w47634 ^ w47632;
	assign w25420 = w47633 ^ w47634;
	assign w6610 = w6734 ^ w6712;
	assign w6609 = w6610 ^ w6611;
	assign w48527 = ~w6609;
	assign w47619 = w48527 ^ w1995;
	assign w20619 = w47619 ^ w47617;
	assign w20621 = w47618 ^ w20619;
	assign w20697 = w47614 ^ w20621;
	assign w20694 = w47615 ^ w20621;
	assign w20696 = w20626 ^ w20621;
	assign w20702 = w47619 ^ w20706;
	assign w20636 = w47619 ^ w47618;
	assign w20689 = w20706 & w20702;
	assign w6604 = w6575 ^ w45485;
	assign w6593 = w45485 ^ w20847;
	assign w48536 = w6592 ^ w6593;
	assign w47610 = w48536 ^ w2004;
	assign w28676 = w47611 ^ w47610;
	assign w28741 = w28676 ^ w28743;
	assign w28747 = w47605 ^ w47610;
	assign w6602 = w6603 ^ w6604;
	assign w48511 = ~w6602;
	assign w47635 = w48511 ^ w1979;
	assign w25443 = w47635 ^ w47633;
	assign w25445 = w47634 ^ w25443;
	assign w25521 = w47630 ^ w25445;
	assign w25518 = w47631 ^ w25445;
	assign w25520 = w25450 ^ w25445;
	assign w25526 = w47635 ^ w25530;
	assign w25460 = w47635 ^ w47634;
	assign w25513 = w25530 & w25526;
	assign w45755 = ~w32503;
	assign w6644 = w32504 ^ w45755;
	assign w6700 = w45755 ^ w45742;
	assign w6634 = w6700 ^ w48705;
	assign w6658 = w6700 ^ w6688;
	assign w45756 = ~w32505;
	assign w6474 = w6683 ^ w45756;
	assign w45757 = ~w32506;
	assign w6431 = w6677 ^ w45757;
	assign w45902 = ~w6030;
	assign w6128 = w45902 ^ w45572;
	assign w6130 = w6129 ^ w6128;
	assign w48350 = ~w6130;
	assign w6132 = w45902 ^ w48458;
	assign w48352 = w6133 ^ w6132;
	assign w6135 = w45902 ^ w48459;
	assign w48353 = w6136 ^ w6135;
	assign w47723 = w48350 ^ w41;
	assign w35978 = w47723 ^ w35982;
	assign w35912 = w47723 ^ w47722;
	assign w35977 = w35912 ^ w35979;
	assign w35985 = w47717 ^ w47723;
	assign w35965 = w35982 & w35978;
	assign w47721 = w48352 ^ w43;
	assign w35895 = w47723 ^ w47721;
	assign w35897 = w47722 ^ w35895;
	assign w35973 = w47718 ^ w35897;
	assign w35970 = w47719 ^ w35897;
	assign w35972 = w35902 ^ w35897;
	assign w35872 = w47721 ^ w47722;
	assign w35966 = w35985 & w35970;
	assign w35900 = w35966 ^ w35896;
	assign w35964 = w35979 & w35972;
	assign w47720 = w48353 ^ w44;
	assign w35898 = w47720 ^ w47718;
	assign w35984 = w47720 ^ w47717;
	assign w35980 = w35984 ^ w35912;
	assign w35976 = w35895 ^ w35984;
	assign w35975 = w47724 ^ w35976;
	assign w35986 = w47722 ^ w47720;
	assign w35971 = w35896 ^ w35986;
	assign w35858 = w35898 ^ w35896;
	assign w35974 = w35895 ^ w35858;
	assign w35857 = w35898 ^ w47719;
	assign w35981 = w47724 ^ w35857;
	assign w35969 = w35976 & w35980;
	assign w35901 = w35969 ^ w35898;
	assign w35968 = w35977 & w35975;
	assign w35967 = w47724 & w35981;
	assign w35963 = w35984 & w35973;
	assign w35899 = w35963 ^ w35897;
	assign w35905 = w35901 ^ w35899;
	assign w35910 = w47717 ^ w35905;
	assign w35962 = w35986 & w35971;
	assign w35919 = w35962 ^ w35968;
	assign w35960 = w35919 ^ w35910;
	assign w35871 = w35962 ^ w35963;
	assign w35918 = w35871 ^ w35872;
	assign w35917 = w35918 ^ w35900;
	assign w35959 = w35965 ^ w35917;
	assign w35961 = w35983 & w35974;
	assign w35956 = w35960 & w35959;
	assign w44874 = w35961 ^ w35964;
	assign w35874 = w35900 ^ w44874;
	assign w35958 = w35874 ^ w35899;
	assign w35955 = w35956 ^ w35958;
	assign w35914 = w35962 ^ w44874;
	assign w35870 = w35965 ^ w35914;
	assign w35952 = w47723 ^ w35870;
	assign w44877 = w35961 ^ w35967;
	assign w35873 = w35905 ^ w44877;
	assign w35916 = w47719 ^ w35873;
	assign w35951 = w35956 ^ w35916;
	assign w35950 = w35951 & w35952;
	assign w35948 = w35956 ^ w35950;
	assign w35869 = w35950 ^ w35914;
	assign w35868 = w35950 ^ w35967;
	assign w35863 = w35868 ^ w35964;
	assign w35947 = w35958 & w35948;
	assign w35945 = w35947 ^ w35955;
	assign w44876 = w35947 ^ w35965;
	assign w35939 = w44876 ^ w35917;
	assign w35928 = w35939 & w35980;
	assign w35937 = w35939 & w35976;
	assign w35906 = w47723 ^ w44876;
	assign w35946 = w35906 ^ w35869;
	assign w35936 = w35946 & w35975;
	assign w35927 = w35946 & w35977;
	assign w35949 = w35950 ^ w35958;
	assign w35935 = w35949 & w47724;
	assign w35926 = w35949 & w35981;
	assign w35911 = w44877 ^ w35896;
	assign w35957 = w35919 ^ w35911;
	assign w35954 = w35957 & w35955;
	assign w35953 = w35954 ^ w35916;
	assign w35865 = w35954 ^ w35966;
	assign w35861 = w35865 ^ w35901;
	assign w35864 = w47717 ^ w35861;
	assign w35941 = w35863 ^ w35864;
	assign w35862 = w35954 ^ w35910;
	assign w35860 = w47719 ^ w35861;
	assign w35944 = w35953 & w35945;
	assign w35909 = w35944 ^ w35919;
	assign w35943 = w35909 ^ w35911;
	assign w35867 = w35944 ^ w35968;
	assign w35859 = w35906 ^ w35867;
	assign w35866 = w35896 ^ w35859;
	assign w35942 = w35863 ^ w35866;
	assign w35940 = w35909 ^ w35862;
	assign w35938 = w35859 ^ w35860;
	assign w35934 = w35940 & w35970;
	assign w35933 = w35943 & w35982;
	assign w35932 = w35953 & w35972;
	assign w35876 = w35932 ^ w35933;
	assign w35931 = w35941 & w35973;
	assign w35930 = w35938 & w35971;
	assign w35891 = w35930 ^ w35933;
	assign w35888 = ~w35891;
	assign w35887 = w35930 ^ w35931;
	assign w35929 = w35942 & w35974;
	assign w35925 = w35940 & w35985;
	assign w35907 = w35925 ^ w35929;
	assign w35892 = w35934 ^ w35925;
	assign w35885 = ~w35907;
	assign w35924 = w35943 & w35978;
	assign w35894 = w35932 ^ w35924;
	assign w35923 = w35953 & w35979;
	assign w35884 = w35885 ^ w35923;
	assign w35922 = w35941 & w35984;
	assign w35921 = w35938 & w35986;
	assign w35920 = w35942 & w35983;
	assign w35886 = w35931 ^ w35920;
	assign w35882 = ~w35886;
	assign w44875 = w35921 ^ w35922;
	assign w35903 = w35927 ^ w44875;
	assign w35904 = w35928 ^ w35903;
	assign w35908 = w35936 ^ w35904;
	assign w35877 = w35935 ^ w35908;
	assign w48700 = w35876 ^ w35877;
	assign w6685 = w48700 ^ w48704;
	assign w6624 = w6685 ^ w6683;
	assign w6470 = w48700 ^ w6471;
	assign w48609 = w6753 ^ w6685;
	assign w47537 = w48609 ^ w1886;
	assign w35913 = w35937 ^ w35908;
	assign w35988 = w35913 ^ w35887;
	assign w35890 = w35894 ^ w44875;
	assign w35889 = w35885 ^ w35890;
	assign w35989 = w35888 ^ w35889;
	assign w44878 = w35933 ^ w35934;
	assign w48701 = w44878 ^ w35913;
	assign w6731 = w48696 ^ w48701;
	assign w6636 = w6731 ^ w6685;
	assign w48634 = w6737 ^ w6731;
	assign w47512 = w48634 ^ w1910;
	assign w6663 = w6677 ^ w48701;
	assign w48610 = w6662 ^ w6663;
	assign w47536 = w48610 ^ w1887;
	assign w6647 = w6731 ^ w6700;
	assign w48619 = w45562 ^ w6647;
	assign w47527 = w48619 ^ w1896;
	assign w35915 = w35930 ^ w44878;
	assign w35881 = w35926 ^ w35915;
	assign w35878 = ~w35881;
	assign w35875 = w35931 ^ w35915;
	assign w48702 = w35904 ^ w35875;
	assign w6666 = w48698 ^ w48702;
	assign w6655 = w6715 ^ w6666;
	assign w48614 = w45757 ^ w6655;
	assign w47532 = w48614 ^ w1891;
	assign w6631 = w6666 ^ w48710;
	assign w6657 = w48702 ^ w32504;
	assign w6619 = w6688 ^ w6666;
	assign w48637 = w48706 ^ w6619;
	assign w47509 = w48637 ^ w1913;
	assign w28614 = w47512 ^ w47509;
	assign w6680 = w48702 ^ w48706;
	assign w6637 = w6680 ^ w48709;
	assign w6761 = ~w6666;
	assign w6654 = w6761 ^ w45756;
	assign w6649 = w6761 ^ w48704;
	assign w6469 = w6761 ^ w48695;
	assign w6738 = w6469 ^ w6470;
	assign w6417 = w6680 ^ w45744;
	assign w6419 = w6680 ^ w48703;
	assign w48618 = w6738 ^ w6682;
	assign w47528 = w48618 ^ w1895;
	assign w44879 = w35935 ^ w35937;
	assign w35893 = w44879 ^ w35890;
	assign w35990 = w35892 ^ w35893;
	assign w35880 = w35884 ^ w44879;
	assign w35883 = w35922 ^ w35880;
	assign w35987 = w35882 ^ w35883;
	assign w35879 = w35903 ^ w35880;
	assign w48699 = w35878 ^ w35879;
	assign w6475 = w45744 ^ w48699;
	assign w48608 = w6474 ^ w6475;
	assign w47538 = w48608 ^ w1885;
	assign w6777 = w47537 ^ w47538;
	assign w6891 = w47538 ^ w47536;
	assign w6705 = w48694 ^ w48699;
	assign w6626 = w6705 ^ w6695;
	assign w48632 = w48703 ^ w6626;
	assign w47514 = w48632 ^ w1908;
	assign w28616 = w47514 ^ w47512;
	assign w28613 = w47509 ^ w47514;
	assign w6420 = w48700 ^ w48699;
	assign w6759 = w6419 ^ w6420;
	assign w48625 = w6759 ^ w6691;
	assign w47521 = w48625 ^ w1902;
	assign w6650 = w6705 ^ w6691;
	assign w6648 = ~w6650;
	assign w48617 = w6648 ^ w6649;
	assign w47529 = w48617 ^ w1894;
	assign w6638 = w6705 ^ w48707;
	assign w48626 = w6636 ^ w6637;
	assign w47520 = w48626 ^ w1903;
	assign w45794 = ~w35988;
	assign w48612 = w45794 ^ w6658;
	assign w6632 = w45563 ^ w45794;
	assign w48629 = w6631 ^ w6632;
	assign w47517 = w48629 ^ w1906;
	assign w20172 = w47520 ^ w47517;
	assign w6730 = w48697 ^ w45794;
	assign w6641 = w6730 ^ w6665;
	assign w48621 = w48698 ^ w6641;
	assign w47525 = w48621 ^ w1898;
	assign w13652 = w47527 ^ w47525;
	assign w13740 = w47528 ^ w47525;
	assign w6620 = w6730 ^ w45742;
	assign w48636 = w6620 ^ w6621;
	assign w47534 = w48612 ^ w1889;
	assign w6803 = w47536 ^ w47534;
	assign w47510 = w48636 ^ w1912;
	assign w28528 = w47512 ^ w47510;
	assign w45795 = ~w35989;
	assign w6639 = w45564 ^ w45795;
	assign w48624 = w6638 ^ w6639;
	assign w47522 = w48624 ^ w1901;
	assign w20174 = w47522 ^ w47520;
	assign w20060 = w47521 ^ w47522;
	assign w20171 = w47517 ^ w47522;
	assign w6432 = w45745 ^ w45795;
	assign w6754 = w6431 ^ w6432;
	assign w48607 = w6754 ^ w6695;
	assign w47539 = w48607 ^ w1884;
	assign w6800 = w47539 ^ w47537;
	assign w6817 = w47539 ^ w47538;
	assign w6802 = w47538 ^ w6800;
	assign w6878 = w47534 ^ w6802;
	assign w6720 = w45756 ^ w45795;
	assign w6651 = w6720 ^ w6683;
	assign w48616 = w48694 ^ w6651;
	assign w6629 = ~w6720;
	assign w6627 = w6629 ^ w6715;
	assign w47530 = w48616 ^ w1893;
	assign w13742 = w47530 ^ w47528;
	assign w13727 = w13652 ^ w13742;
	assign w13628 = w47529 ^ w47530;
	assign w13739 = w47525 ^ w47530;
	assign w13718 = w13742 & w13727;
	assign w45796 = ~w35990;
	assign w6728 = w45757 ^ w45796;
	assign w6653 = w6728 ^ w6695;
	assign w6652 = w6653 ^ w6654;
	assign w6630 = w6728 ^ w6665;
	assign w48630 = w45565 ^ w6630;
	assign w47516 = w48630 ^ w45167;
	assign w28532 = w47516 ^ w47510;
	assign w48615 = ~w6652;
	assign w47531 = w48615 ^ w1892;
	assign w13651 = w47531 ^ w47529;
	assign w13653 = w47530 ^ w13651;
	assign w13726 = w47527 ^ w13653;
	assign w13732 = w13651 ^ w13740;
	assign w13731 = w47532 ^ w13732;
	assign w13668 = w47531 ^ w47530;
	assign w13736 = w13740 ^ w13668;
	assign w13741 = w47525 ^ w47531;
	assign w13725 = w13732 & w13736;
	assign w13722 = w13741 & w13726;
	assign w13656 = w13722 ^ w13652;
	assign w6640 = w6728 ^ w6680;
	assign w48622 = w45745 ^ w6640;
	assign w48606 = w45796 ^ w6476;
	assign w47540 = w48606 ^ w1883;
	assign w6807 = w47540 ^ w47534;
	assign w6877 = w6807 ^ w6802;
	assign w47524 = w48622 ^ w1899;
	assign w6418 = w45565 ^ w45796;
	assign w6760 = w6417 ^ w6418;
	assign w48623 = w6760 ^ w6720;
	assign w47523 = w48623 ^ w1900;
	assign w20083 = w47523 ^ w47521;
	assign w20085 = w47522 ^ w20083;
	assign w20164 = w20083 ^ w20172;
	assign w20163 = w47524 ^ w20164;
	assign w20100 = w47523 ^ w47522;
	assign w20168 = w20172 ^ w20100;
	assign w20173 = w47517 ^ w47523;
	assign w20157 = w20164 & w20168;
	assign w45801 = ~w35987;
	assign w6690 = w45801 ^ w45562;
	assign w6633 = w6730 ^ w6690;
	assign w6635 = w45801 ^ w48701;
	assign w6643 = w6688 ^ w45801;
	assign w6642 = w6643 ^ w6644;
	assign w6661 = ~w6690;
	assign w6659 = w6661 ^ w45742;
	assign w48611 = w6659 ^ w6660;
	assign w47535 = w48611 ^ w1888;
	assign w48628 = w45743 ^ w6633;
	assign w47518 = w48628 ^ w1905;
	assign w20161 = w47518 ^ w20085;
	assign w20086 = w47520 ^ w47518;
	assign w20089 = w20157 ^ w20086;
	assign w20090 = w47524 ^ w47518;
	assign w20160 = w20090 ^ w20085;
	assign w20151 = w20172 & w20161;
	assign w20087 = w20151 ^ w20085;
	assign w20093 = w20089 ^ w20087;
	assign w20098 = w47517 ^ w20093;
	assign w48627 = w6634 ^ w6635;
	assign w47519 = w48627 ^ w1904;
	assign w20158 = w47519 ^ w20085;
	assign w20084 = w47519 ^ w47517;
	assign w20159 = w20084 ^ w20174;
	assign w20167 = w20084 ^ w20090;
	assign w20165 = w20100 ^ w20167;
	assign w20170 = w47519 ^ w20090;
	assign w20166 = w47523 ^ w20170;
	assign w20046 = w20086 ^ w20084;
	assign w20162 = w20083 ^ w20046;
	assign w20045 = w20086 ^ w47519;
	assign w20169 = w47524 ^ w20045;
	assign w20156 = w20165 & w20163;
	assign w20155 = w47524 & w20169;
	assign w20154 = w20173 & w20158;
	assign w20088 = w20154 ^ w20084;
	assign w20153 = w20170 & w20166;
	assign w20152 = w20167 & w20160;
	assign w20150 = w20174 & w20159;
	assign w20107 = w20150 ^ w20156;
	assign w20148 = w20107 ^ w20098;
	assign w20059 = w20150 ^ w20151;
	assign w20106 = w20059 ^ w20060;
	assign w20105 = w20106 ^ w20088;
	assign w20147 = w20153 ^ w20105;
	assign w20149 = w20171 & w20162;
	assign w20144 = w20148 & w20147;
	assign w48620 = ~w6642;
	assign w47526 = w48620 ^ w1897;
	assign w13729 = w47526 ^ w13653;
	assign w13654 = w47528 ^ w47526;
	assign w13657 = w13725 ^ w13654;
	assign w13658 = w47532 ^ w47526;
	assign w13728 = w13658 ^ w13653;
	assign w13735 = w13652 ^ w13658;
	assign w13733 = w13668 ^ w13735;
	assign w13738 = w47527 ^ w13658;
	assign w13734 = w47531 ^ w13738;
	assign w13614 = w13654 ^ w13652;
	assign w13730 = w13651 ^ w13614;
	assign w13613 = w13654 ^ w47527;
	assign w13737 = w47532 ^ w13613;
	assign w13724 = w13733 & w13731;
	assign w13675 = w13718 ^ w13724;
	assign w13723 = w47532 & w13737;
	assign w13721 = w13738 & w13734;
	assign w13720 = w13735 & w13728;
	assign w13719 = w13740 & w13729;
	assign w13655 = w13719 ^ w13653;
	assign w13661 = w13657 ^ w13655;
	assign w13666 = w47525 ^ w13661;
	assign w13716 = w13675 ^ w13666;
	assign w13627 = w13718 ^ w13719;
	assign w13674 = w13627 ^ w13628;
	assign w13673 = w13674 ^ w13656;
	assign w13715 = w13721 ^ w13673;
	assign w13717 = w13739 & w13730;
	assign w13712 = w13716 & w13715;
	assign w6622 = w6690 ^ w6682;
	assign w48635 = w45755 ^ w6622;
	assign w47511 = w48635 ^ w1911;
	assign w28526 = w47511 ^ w47509;
	assign w28601 = w28526 ^ w28616;
	assign w28609 = w28526 ^ w28532;
	assign w28612 = w47511 ^ w28532;
	assign w28488 = w28528 ^ w28526;
	assign w28487 = w28528 ^ w47511;
	assign w28611 = w47516 ^ w28487;
	assign w28597 = w47516 & w28611;
	assign w28592 = w28616 & w28601;
	assign w6887 = w47535 ^ w6807;
	assign w6883 = w47539 ^ w6887;
	assign w6762 = w6803 ^ w47535;
	assign w6886 = w47540 ^ w6762;
	assign w6872 = w47540 & w6886;
	assign w6870 = w6887 & w6883;
	assign w43942 = w13717 ^ w13723;
	assign w13667 = w43942 ^ w13652;
	assign w13713 = w13675 ^ w13667;
	assign w13629 = w13661 ^ w43942;
	assign w13672 = w47527 ^ w13629;
	assign w13707 = w13712 ^ w13672;
	assign w43943 = w13717 ^ w13720;
	assign w13670 = w13718 ^ w43943;
	assign w13626 = w13721 ^ w13670;
	assign w13708 = w47531 ^ w13626;
	assign w13706 = w13707 & w13708;
	assign w13704 = w13712 ^ w13706;
	assign w13625 = w13706 ^ w13670;
	assign w13624 = w13706 ^ w13723;
	assign w13619 = w13624 ^ w13720;
	assign w13630 = w13656 ^ w43943;
	assign w13714 = w13630 ^ w13655;
	assign w13705 = w13706 ^ w13714;
	assign w13711 = w13712 ^ w13714;
	assign w13710 = w13713 & w13711;
	assign w13709 = w13710 ^ w13672;
	assign w13621 = w13710 ^ w13722;
	assign w13617 = w13621 ^ w13657;
	assign w13620 = w47525 ^ w13617;
	assign w13697 = w13619 ^ w13620;
	assign w13618 = w13710 ^ w13666;
	assign w13616 = w47527 ^ w13617;
	assign w13703 = w13714 & w13704;
	assign w13701 = w13703 ^ w13711;
	assign w13700 = w13709 & w13701;
	assign w13665 = w13700 ^ w13675;
	assign w13699 = w13665 ^ w13667;
	assign w13623 = w13700 ^ w13724;
	assign w13696 = w13665 ^ w13618;
	assign w13691 = w13705 & w47532;
	assign w13690 = w13696 & w13726;
	assign w13689 = w13699 & w13738;
	assign w13688 = w13709 & w13728;
	assign w13632 = w13688 ^ w13689;
	assign w13687 = w13697 & w13729;
	assign w13682 = w13705 & w13737;
	assign w13681 = w13696 & w13741;
	assign w13648 = w13690 ^ w13681;
	assign w13680 = w13699 & w13734;
	assign w13650 = w13688 ^ w13680;
	assign w13679 = w13709 & w13735;
	assign w13678 = w13697 & w13740;
	assign w43944 = w13689 ^ w13690;
	assign w43946 = w13703 ^ w13721;
	assign w13662 = w47531 ^ w43946;
	assign w13615 = w13662 ^ w13623;
	assign w13622 = w13652 ^ w13615;
	assign w13698 = w13619 ^ w13622;
	assign w13685 = w13698 & w13730;
	assign w13663 = w13681 ^ w13685;
	assign w13641 = ~w13663;
	assign w13694 = w13615 ^ w13616;
	assign w13686 = w13694 & w13727;
	assign w13643 = w13686 ^ w13687;
	assign w13671 = w13686 ^ w43944;
	assign w13637 = w13682 ^ w13671;
	assign w13634 = ~w13637;
	assign w13631 = w13687 ^ w13671;
	assign w13647 = w13686 ^ w13689;
	assign w13644 = ~w13647;
	assign w13640 = w13641 ^ w13679;
	assign w13677 = w13694 & w13742;
	assign w13676 = w13698 & w13739;
	assign w13642 = w13687 ^ w13676;
	assign w13638 = ~w13642;
	assign w43535 = w13677 ^ w13678;
	assign w13646 = w13650 ^ w43535;
	assign w13645 = w13641 ^ w13646;
	assign w13745 = w13644 ^ w13645;
	assign w48863 = ~w13745;
	assign w13702 = w13662 ^ w13625;
	assign w13683 = w13702 & w13733;
	assign w13692 = w13702 & w13731;
	assign w13659 = w13683 ^ w43535;
	assign w13695 = w43946 ^ w13673;
	assign w13693 = w13695 & w13732;
	assign w13684 = w13695 & w13736;
	assign w13660 = w13684 ^ w13659;
	assign w13664 = w13692 ^ w13660;
	assign w13669 = w13693 ^ w13664;
	assign w48866 = w43944 ^ w13669;
	assign w13744 = w13669 ^ w13643;
	assign w13633 = w13691 ^ w13664;
	assign w48865 = w13632 ^ w13633;
	assign w48867 = w13660 ^ w13631;
	assign w6907 = ~w48865;
	assign w43945 = w13691 ^ w13693;
	assign w13649 = w43945 ^ w13646;
	assign w13746 = w13648 ^ w13649;
	assign w13636 = w13640 ^ w43945;
	assign w13639 = w13678 ^ w13636;
	assign w13743 = w13638 ^ w13639;
	assign w13635 = w13659 ^ w13636;
	assign w48864 = w13634 ^ w13635;
	assign w44210 = w20149 ^ w20152;
	assign w20062 = w20088 ^ w44210;
	assign w20146 = w20062 ^ w20087;
	assign w20143 = w20144 ^ w20146;
	assign w20102 = w20150 ^ w44210;
	assign w20058 = w20153 ^ w20102;
	assign w20140 = w47523 ^ w20058;
	assign w44213 = w20149 ^ w20155;
	assign w20061 = w20093 ^ w44213;
	assign w20104 = w47519 ^ w20061;
	assign w20139 = w20144 ^ w20104;
	assign w20138 = w20139 & w20140;
	assign w20136 = w20144 ^ w20138;
	assign w20057 = w20138 ^ w20102;
	assign w20056 = w20138 ^ w20155;
	assign w20051 = w20056 ^ w20152;
	assign w20135 = w20146 & w20136;
	assign w20133 = w20135 ^ w20143;
	assign w44212 = w20135 ^ w20153;
	assign w20127 = w44212 ^ w20105;
	assign w20116 = w20127 & w20168;
	assign w20125 = w20127 & w20164;
	assign w20094 = w47523 ^ w44212;
	assign w20134 = w20094 ^ w20057;
	assign w20124 = w20134 & w20163;
	assign w20115 = w20134 & w20165;
	assign w20137 = w20138 ^ w20146;
	assign w20123 = w20137 & w47524;
	assign w20114 = w20137 & w20169;
	assign w20099 = w44213 ^ w20084;
	assign w20145 = w20107 ^ w20099;
	assign w20142 = w20145 & w20143;
	assign w20141 = w20142 ^ w20104;
	assign w20053 = w20142 ^ w20154;
	assign w20049 = w20053 ^ w20089;
	assign w20052 = w47517 ^ w20049;
	assign w20129 = w20051 ^ w20052;
	assign w20050 = w20142 ^ w20098;
	assign w20048 = w47519 ^ w20049;
	assign w20132 = w20141 & w20133;
	assign w20097 = w20132 ^ w20107;
	assign w20131 = w20097 ^ w20099;
	assign w20055 = w20132 ^ w20156;
	assign w20047 = w20094 ^ w20055;
	assign w20054 = w20084 ^ w20047;
	assign w20130 = w20051 ^ w20054;
	assign w20128 = w20097 ^ w20050;
	assign w20126 = w20047 ^ w20048;
	assign w20122 = w20128 & w20158;
	assign w20121 = w20131 & w20170;
	assign w20120 = w20141 & w20160;
	assign w20064 = w20120 ^ w20121;
	assign w20119 = w20129 & w20161;
	assign w20118 = w20126 & w20159;
	assign w20079 = w20118 ^ w20121;
	assign w20076 = ~w20079;
	assign w20075 = w20118 ^ w20119;
	assign w20117 = w20130 & w20162;
	assign w20113 = w20128 & w20173;
	assign w20095 = w20113 ^ w20117;
	assign w20080 = w20122 ^ w20113;
	assign w20073 = ~w20095;
	assign w20112 = w20131 & w20166;
	assign w20082 = w20120 ^ w20112;
	assign w20111 = w20141 & w20167;
	assign w20072 = w20073 ^ w20111;
	assign w20110 = w20129 & w20172;
	assign w20109 = w20126 & w20174;
	assign w20108 = w20130 & w20171;
	assign w20074 = w20119 ^ w20108;
	assign w20070 = ~w20074;
	assign w44211 = w20109 ^ w20110;
	assign w20091 = w20115 ^ w44211;
	assign w20092 = w20116 ^ w20091;
	assign w20096 = w20124 ^ w20092;
	assign w20065 = w20123 ^ w20096;
	assign w48851 = w20064 ^ w20065;
	assign w20101 = w20125 ^ w20096;
	assign w20176 = w20101 ^ w20075;
	assign w20078 = w20082 ^ w44211;
	assign w20077 = w20073 ^ w20078;
	assign w20177 = w20076 ^ w20077;
	assign w48849 = ~w20177;
	assign w44214 = w20121 ^ w20122;
	assign w48852 = w44214 ^ w20101;
	assign w20103 = w20118 ^ w44214;
	assign w20069 = w20114 ^ w20103;
	assign w20066 = ~w20069;
	assign w20063 = w20119 ^ w20103;
	assign w48853 = w20092 ^ w20063;
	assign w44215 = w20123 ^ w20125;
	assign w20081 = w44215 ^ w20078;
	assign w20178 = w20080 ^ w20081;
	assign w20068 = w20072 ^ w44215;
	assign w20071 = w20110 ^ w20068;
	assign w20175 = w20070 ^ w20071;
	assign w20067 = w20091 ^ w20068;
	assign w48850 = w20066 ^ w20067;
	assign w6947 = ~w48850;
	assign w6946 = w48851 ^ w6947;
	assign w6875 = w47535 ^ w6802;
	assign w45271 = ~w13743;
	assign w45272 = ~w13744;
	assign w7030 = w45272 ^ w45271;
	assign w45273 = ~w13746;
	assign w45446 = ~w20175;
	assign w45447 = ~w20176;
	assign w45448 = ~w20178;
	assign w45903 = ~w6032;
	assign w6210 = w45903 ^ w45494;
	assign w48398 = w6211 ^ w6210;
	assign w6218 = w45903 ^ w48487;
	assign w48401 = w6219 ^ w6218;
	assign w6215 = w45903 ^ w48486;
	assign w48400 = w6216 ^ w6215;
	assign w47673 = w48400 ^ w91;
	assign w32120 = w47673 ^ w47674;
	assign w47675 = w48398 ^ w89;
	assign w32143 = w47675 ^ w47673;
	assign w32145 = w47674 ^ w32143;
	assign w32221 = w47670 ^ w32145;
	assign w32218 = w47671 ^ w32145;
	assign w32220 = w32150 ^ w32145;
	assign w32226 = w47675 ^ w32230;
	assign w32160 = w47675 ^ w47674;
	assign w32225 = w32160 ^ w32227;
	assign w32233 = w47669 ^ w47675;
	assign w32214 = w32233 & w32218;
	assign w32148 = w32214 ^ w32144;
	assign w32213 = w32230 & w32226;
	assign w32212 = w32227 & w32220;
	assign w47672 = w48401 ^ w92;
	assign w32146 = w47672 ^ w47670;
	assign w32232 = w47672 ^ w47669;
	assign w32228 = w32232 ^ w32160;
	assign w32224 = w32143 ^ w32232;
	assign w32223 = w47676 ^ w32224;
	assign w32234 = w47674 ^ w47672;
	assign w32219 = w32144 ^ w32234;
	assign w32106 = w32146 ^ w32144;
	assign w32222 = w32143 ^ w32106;
	assign w32105 = w32146 ^ w47671;
	assign w32229 = w47676 ^ w32105;
	assign w32217 = w32224 & w32228;
	assign w32149 = w32217 ^ w32146;
	assign w32216 = w32225 & w32223;
	assign w32215 = w47676 & w32229;
	assign w32211 = w32232 & w32221;
	assign w32147 = w32211 ^ w32145;
	assign w32153 = w32149 ^ w32147;
	assign w32158 = w47669 ^ w32153;
	assign w32210 = w32234 & w32219;
	assign w32167 = w32210 ^ w32216;
	assign w32208 = w32167 ^ w32158;
	assign w32119 = w32210 ^ w32211;
	assign w32166 = w32119 ^ w32120;
	assign w32165 = w32166 ^ w32148;
	assign w32207 = w32213 ^ w32165;
	assign w32209 = w32231 & w32222;
	assign w32204 = w32208 & w32207;
	assign w44717 = w32209 ^ w32215;
	assign w32159 = w44717 ^ w32144;
	assign w32205 = w32167 ^ w32159;
	assign w32121 = w32153 ^ w44717;
	assign w32164 = w47671 ^ w32121;
	assign w32199 = w32204 ^ w32164;
	assign w44718 = w32209 ^ w32212;
	assign w32162 = w32210 ^ w44718;
	assign w32118 = w32213 ^ w32162;
	assign w32200 = w47675 ^ w32118;
	assign w32198 = w32199 & w32200;
	assign w32117 = w32198 ^ w32162;
	assign w32116 = w32198 ^ w32215;
	assign w32111 = w32116 ^ w32212;
	assign w32196 = w32204 ^ w32198;
	assign w32122 = w32148 ^ w44718;
	assign w32206 = w32122 ^ w32147;
	assign w32197 = w32198 ^ w32206;
	assign w32203 = w32204 ^ w32206;
	assign w32202 = w32205 & w32203;
	assign w32201 = w32202 ^ w32164;
	assign w32113 = w32202 ^ w32214;
	assign w32109 = w32113 ^ w32149;
	assign w32112 = w47669 ^ w32109;
	assign w32189 = w32111 ^ w32112;
	assign w32110 = w32202 ^ w32158;
	assign w32108 = w47671 ^ w32109;
	assign w32195 = w32206 & w32196;
	assign w32193 = w32195 ^ w32203;
	assign w32192 = w32201 & w32193;
	assign w32157 = w32192 ^ w32167;
	assign w32191 = w32157 ^ w32159;
	assign w32115 = w32192 ^ w32216;
	assign w32188 = w32157 ^ w32110;
	assign w32183 = w32197 & w47676;
	assign w32182 = w32188 & w32218;
	assign w32181 = w32191 & w32230;
	assign w32180 = w32201 & w32220;
	assign w32124 = w32180 ^ w32181;
	assign w32179 = w32189 & w32221;
	assign w32174 = w32197 & w32229;
	assign w32173 = w32188 & w32233;
	assign w32140 = w32182 ^ w32173;
	assign w32172 = w32191 & w32226;
	assign w32142 = w32180 ^ w32172;
	assign w32171 = w32201 & w32227;
	assign w32170 = w32189 & w32232;
	assign w44719 = w32181 ^ w32182;
	assign w44721 = w32195 ^ w32213;
	assign w32154 = w47675 ^ w44721;
	assign w32194 = w32154 ^ w32117;
	assign w32175 = w32194 & w32225;
	assign w32184 = w32194 & w32223;
	assign w32107 = w32154 ^ w32115;
	assign w32114 = w32144 ^ w32107;
	assign w32190 = w32111 ^ w32114;
	assign w32177 = w32190 & w32222;
	assign w32155 = w32173 ^ w32177;
	assign w32133 = ~w32155;
	assign w32132 = w32133 ^ w32171;
	assign w32186 = w32107 ^ w32108;
	assign w32169 = w32186 & w32234;
	assign w32168 = w32190 & w32231;
	assign w32134 = w32179 ^ w32168;
	assign w32130 = ~w32134;
	assign w43588 = w32169 ^ w32170;
	assign w32151 = w32175 ^ w43588;
	assign w32138 = w32142 ^ w43588;
	assign w32137 = w32133 ^ w32138;
	assign w32178 = w32186 & w32219;
	assign w32139 = w32178 ^ w32181;
	assign w32136 = ~w32139;
	assign w32237 = w32136 ^ w32137;
	assign w32135 = w32178 ^ w32179;
	assign w32163 = w32178 ^ w44719;
	assign w32123 = w32179 ^ w32163;
	assign w32129 = w32174 ^ w32163;
	assign w32126 = ~w32129;
	assign w32187 = w44721 ^ w32165;
	assign w32185 = w32187 & w32224;
	assign w32176 = w32187 & w32228;
	assign w32152 = w32176 ^ w32151;
	assign w32156 = w32184 ^ w32152;
	assign w32161 = w32185 ^ w32156;
	assign w48692 = w44719 ^ w32161;
	assign w32236 = w32161 ^ w32135;
	assign w32125 = w32183 ^ w32156;
	assign w48691 = w32124 ^ w32125;
	assign w48693 = w32152 ^ w32123;
	assign w6675 = w48678 ^ w48693;
	assign w6707 = w48687 ^ w48691;
	assign w6698 = w48688 ^ w48692;
	assign w6456 = w6455 ^ w48692;
	assign w6744 = w6456 ^ w6457;
	assign w48594 = w6744 ^ w6710;
	assign w6452 = w6455 ^ w48691;
	assign w6745 = w6452 ^ w6453;
	assign w48593 = w6745 ^ w6718;
	assign w47553 = w48593 ^ w1933;
	assign w6510 = w6501 ^ w6707;
	assign w48585 = w6510 ^ w6511;
	assign w47561 = w48585 ^ w1925;
	assign w6667 = w48689 ^ w48693;
	assign w6508 = w6485 ^ w6698;
	assign w6505 = w6696 ^ w6667;
	assign w48586 = w6508 ^ w6509;
	assign w6492 = w45888 ^ w48693;
	assign w6491 = w6733 ^ w6667;
	assign w48598 = w45474 ^ w6491;
	assign w47548 = w48598 ^ w1938;
	assign w48589 = w48678 ^ w6505;
	assign w48597 = w6492 ^ w6493;
	assign w47549 = w48597 ^ w1937;
	assign w6480 = w6482 ^ w6707;
	assign w6479 = w6703 ^ w6698;
	assign w48603 = w45479 ^ w6479;
	assign w47543 = w48603 ^ w1943;
	assign w6448 = w6675 ^ w48691;
	assign w6747 = w6448 ^ w6449;
	assign w48578 = w6747 ^ w6698;
	assign w47568 = w48578 ^ w1918;
	assign w47552 = w48594 ^ w1934;
	assign w20306 = w47552 ^ w47549;
	assign w47560 = w48586 ^ w1926;
	assign w6444 = ~w6675;
	assign w47557 = w48589 ^ w1929;
	assign w34376 = w47560 ^ w47557;
	assign w44720 = w32183 ^ w32185;
	assign w32141 = w44720 ^ w32138;
	assign w32238 = w32140 ^ w32141;
	assign w32128 = w32132 ^ w44720;
	assign w32131 = w32170 ^ w32128;
	assign w32235 = w32130 ^ w32131;
	assign w32127 = w32151 ^ w32128;
	assign w48690 = w32126 ^ w32127;
	assign w6717 = w48686 ^ w48690;
	assign w6530 = ~w6717;
	assign w6512 = w6732 ^ w6717;
	assign w48584 = w48675 ^ w6512;
	assign w47562 = w48584 ^ w1924;
	assign w34378 = w47562 ^ w47560;
	assign w34264 = w47561 ^ w47562;
	assign w34375 = w47557 ^ w47562;
	assign w6499 = w6501 ^ w48690;
	assign w48592 = w6499 ^ w6500;
	assign w47554 = w48592 ^ w1932;
	assign w20308 = w47554 ^ w47552;
	assign w20194 = w47553 ^ w47554;
	assign w20305 = w47549 ^ w47554;
	assign w6483 = w6485 ^ w6717;
	assign w6445 = w6444 ^ w48690;
	assign w6748 = w6445 ^ w6446;
	assign w48577 = w6748 ^ w6707;
	assign w47569 = w48577 ^ w1917;
	assign w45746 = ~w32235;
	assign w6497 = w6703 ^ w45746;
	assign w48595 = w6497 ^ w6498;
	assign w47551 = w48595 ^ w1935;
	assign w20218 = w47551 ^ w47549;
	assign w20293 = w20218 ^ w20308;
	assign w20284 = w20308 & w20293;
	assign w6692 = w45479 ^ w45746;
	assign w6478 = w6696 ^ w6692;
	assign w6527 = w6692 ^ w48692;
	assign w6525 = ~w6527;
	assign w48579 = w6525 ^ w6526;
	assign w47567 = w48579 ^ w1919;
	assign w6507 = w6710 ^ w6692;
	assign w48587 = w45471 ^ w6507;
	assign w47559 = w48587 ^ w1927;
	assign w34288 = w47559 ^ w47557;
	assign w34363 = w34288 ^ w34378;
	assign w34354 = w34378 & w34363;
	assign w48604 = w45480 ^ w6478;
	assign w47542 = w48604 ^ w1944;
	assign w31748 = w47548 ^ w47542;
	assign w31828 = w47543 ^ w31748;
	assign w45747 = ~w32236;
	assign w6517 = w6667 ^ w45747;
	assign w48581 = w6517 ^ w6518;
	assign w47565 = w48581 ^ w1921;
	assign w20352 = w47567 ^ w47565;
	assign w20440 = w47568 ^ w47565;
	assign w6496 = w6696 ^ w45747;
	assign w6494 = ~w6496;
	assign w48596 = w6494 ^ w6495;
	assign w47550 = w48596 ^ w1936;
	assign w20220 = w47552 ^ w47550;
	assign w20180 = w20220 ^ w20218;
	assign w20179 = w20220 ^ w47551;
	assign w6681 = w45480 ^ w45747;
	assign w6477 = w6681 ^ w6670;
	assign w48605 = w48689 ^ w6477;
	assign w47541 = w48605 ^ w1945;
	assign w31742 = w47543 ^ w47541;
	assign w31825 = w31742 ^ w31748;
	assign w6520 = w6681 ^ w45746;
	assign w6519 = w6520 ^ w6521;
	assign w48580 = ~w6519;
	assign w47566 = w48580 ^ w1920;
	assign w20354 = w47568 ^ w47566;
	assign w20314 = w20354 ^ w20352;
	assign w20313 = w20354 ^ w47567;
	assign w6506 = w6703 ^ w6681;
	assign w48588 = w45472 ^ w6506;
	assign w47558 = w48588 ^ w1928;
	assign w34290 = w47560 ^ w47558;
	assign w34250 = w34290 ^ w34288;
	assign w34249 = w34290 ^ w47559;
	assign w45748 = ~w32237;
	assign w6721 = w45481 ^ w45748;
	assign w6450 = w6674 ^ w45748;
	assign w6746 = w6450 ^ w6451;
	assign w48591 = w6746 ^ w6732;
	assign w6528 = w6530 ^ w45748;
	assign w48576 = w6528 ^ w6529;
	assign w47570 = w48576 ^ w1916;
	assign w20442 = w47570 ^ w47568;
	assign w20427 = w20352 ^ w20442;
	assign w20328 = w47569 ^ w47570;
	assign w20439 = w47565 ^ w47570;
	assign w20418 = w20442 & w20427;
	assign w6514 = w6733 ^ w6721;
	assign w6513 = w6514 ^ w6515;
	assign w48583 = ~w6513;
	assign w47563 = w48583 ^ w1923;
	assign w34287 = w47563 ^ w47561;
	assign w34289 = w47562 ^ w34287;
	assign w34365 = w47558 ^ w34289;
	assign w34362 = w47559 ^ w34289;
	assign w34368 = w34287 ^ w34376;
	assign w34304 = w47563 ^ w47562;
	assign w34372 = w34376 ^ w34304;
	assign w34366 = w34287 ^ w34250;
	assign w34377 = w47557 ^ w47563;
	assign w34361 = w34368 & w34372;
	assign w34293 = w34361 ^ w34290;
	assign w34358 = w34377 & w34362;
	assign w34292 = w34358 ^ w34288;
	assign w34355 = w34376 & w34365;
	assign w34291 = w34355 ^ w34289;
	assign w34297 = w34293 ^ w34291;
	assign w34302 = w47557 ^ w34297;
	assign w34263 = w34354 ^ w34355;
	assign w34310 = w34263 ^ w34264;
	assign w34309 = w34310 ^ w34292;
	assign w34353 = w34375 & w34366;
	assign w6486 = w6725 ^ w6721;
	assign w48600 = w48686 ^ w6486;
	assign w47546 = w48600 ^ w1940;
	assign w31829 = w47541 ^ w47546;
	assign w47555 = w48591 ^ w1931;
	assign w20217 = w47555 ^ w47553;
	assign w20219 = w47554 ^ w20217;
	assign w20295 = w47550 ^ w20219;
	assign w20292 = w47551 ^ w20219;
	assign w20298 = w20217 ^ w20306;
	assign w20234 = w47555 ^ w47554;
	assign w20302 = w20306 ^ w20234;
	assign w20296 = w20217 ^ w20180;
	assign w20307 = w47549 ^ w47555;
	assign w20291 = w20298 & w20302;
	assign w20223 = w20291 ^ w20220;
	assign w20288 = w20307 & w20292;
	assign w20222 = w20288 ^ w20218;
	assign w20285 = w20306 & w20295;
	assign w20221 = w20285 ^ w20219;
	assign w20227 = w20223 ^ w20221;
	assign w20232 = w47549 ^ w20227;
	assign w20193 = w20284 ^ w20285;
	assign w20240 = w20193 ^ w20194;
	assign w20239 = w20240 ^ w20222;
	assign w20283 = w20305 & w20296;
	assign w45749 = ~w32238;
	assign w6729 = w45474 ^ w45749;
	assign w6531 = w6729 ^ w6675;
	assign w48574 = w45785 ^ w6531;
	assign w6516 = w6729 ^ w6670;
	assign w48582 = w45466 ^ w6516;
	assign w47564 = w48582 ^ w1922;
	assign w34367 = w47564 ^ w34368;
	assign w34294 = w47564 ^ w47558;
	assign w34364 = w34294 ^ w34289;
	assign w34371 = w34288 ^ w34294;
	assign w34369 = w34304 ^ w34371;
	assign w34374 = w47559 ^ w34294;
	assign w34370 = w47563 ^ w34374;
	assign w34373 = w47564 ^ w34249;
	assign w34360 = w34369 & w34367;
	assign w34311 = w34354 ^ w34360;
	assign w34352 = w34311 ^ w34302;
	assign w34359 = w47564 & w34373;
	assign w34357 = w34374 & w34370;
	assign w34351 = w34357 ^ w34309;
	assign w34356 = w34371 & w34364;
	assign w34348 = w34352 & w34351;
	assign w48590 = w45749 ^ w6502;
	assign w6490 = w6732 ^ w6729;
	assign w6488 = ~w6490;
	assign w6442 = w6444 ^ w45749;
	assign w6749 = w6442 ^ w6443;
	assign w48575 = w6749 ^ w6721;
	assign w47571 = w48575 ^ w1915;
	assign w20351 = w47571 ^ w47569;
	assign w20353 = w47570 ^ w20351;
	assign w20429 = w47566 ^ w20353;
	assign w20426 = w47567 ^ w20353;
	assign w20432 = w20351 ^ w20440;
	assign w20368 = w47571 ^ w47570;
	assign w20436 = w20440 ^ w20368;
	assign w20430 = w20351 ^ w20314;
	assign w20441 = w47565 ^ w47571;
	assign w20425 = w20432 & w20436;
	assign w20357 = w20425 ^ w20354;
	assign w20422 = w20441 & w20426;
	assign w20356 = w20422 ^ w20352;
	assign w20419 = w20440 & w20429;
	assign w20355 = w20419 ^ w20353;
	assign w20361 = w20357 ^ w20355;
	assign w20366 = w47565 ^ w20361;
	assign w20327 = w20418 ^ w20419;
	assign w20374 = w20327 ^ w20328;
	assign w20373 = w20374 ^ w20356;
	assign w20417 = w20439 & w20430;
	assign w47556 = w48590 ^ w1930;
	assign w20297 = w47556 ^ w20298;
	assign w20224 = w47556 ^ w47550;
	assign w20294 = w20224 ^ w20219;
	assign w20301 = w20218 ^ w20224;
	assign w20299 = w20234 ^ w20301;
	assign w20304 = w47551 ^ w20224;
	assign w20300 = w47555 ^ w20304;
	assign w20303 = w47556 ^ w20179;
	assign w20290 = w20299 & w20297;
	assign w20241 = w20284 ^ w20290;
	assign w20282 = w20241 ^ w20232;
	assign w20289 = w47556 & w20303;
	assign w20287 = w20304 & w20300;
	assign w20281 = w20287 ^ w20239;
	assign w20286 = w20301 & w20294;
	assign w20278 = w20282 & w20281;
	assign w44216 = w20283 ^ w20289;
	assign w20195 = w20227 ^ w44216;
	assign w20238 = w47551 ^ w20195;
	assign w20273 = w20278 ^ w20238;
	assign w20233 = w44216 ^ w20218;
	assign w20279 = w20241 ^ w20233;
	assign w44217 = w20283 ^ w20286;
	assign w20236 = w20284 ^ w44217;
	assign w20192 = w20287 ^ w20236;
	assign w20274 = w47555 ^ w20192;
	assign w20272 = w20273 & w20274;
	assign w20270 = w20278 ^ w20272;
	assign w20191 = w20272 ^ w20236;
	assign w20190 = w20272 ^ w20289;
	assign w20185 = w20190 ^ w20286;
	assign w20196 = w20222 ^ w44217;
	assign w20280 = w20196 ^ w20221;
	assign w20271 = w20272 ^ w20280;
	assign w20277 = w20278 ^ w20280;
	assign w20276 = w20279 & w20277;
	assign w20275 = w20276 ^ w20238;
	assign w20187 = w20276 ^ w20288;
	assign w20183 = w20187 ^ w20223;
	assign w20186 = w47549 ^ w20183;
	assign w20263 = w20185 ^ w20186;
	assign w20184 = w20276 ^ w20232;
	assign w20182 = w47551 ^ w20183;
	assign w20269 = w20280 & w20270;
	assign w20267 = w20269 ^ w20277;
	assign w20266 = w20275 & w20267;
	assign w20231 = w20266 ^ w20241;
	assign w20265 = w20231 ^ w20233;
	assign w20189 = w20266 ^ w20290;
	assign w20262 = w20231 ^ w20184;
	assign w20257 = w20271 & w47556;
	assign w20256 = w20262 & w20292;
	assign w20255 = w20265 & w20304;
	assign w20254 = w20275 & w20294;
	assign w20198 = w20254 ^ w20255;
	assign w20253 = w20263 & w20295;
	assign w20248 = w20271 & w20303;
	assign w20247 = w20262 & w20307;
	assign w20214 = w20256 ^ w20247;
	assign w20246 = w20265 & w20300;
	assign w20216 = w20254 ^ w20246;
	assign w20245 = w20275 & w20301;
	assign w20244 = w20263 & w20306;
	assign w44219 = w20255 ^ w20256;
	assign w44221 = w20269 ^ w20287;
	assign w20261 = w44221 ^ w20239;
	assign w20250 = w20261 & w20302;
	assign w20259 = w20261 & w20298;
	assign w44220 = w20257 ^ w20259;
	assign w20228 = w47555 ^ w44221;
	assign w20268 = w20228 ^ w20191;
	assign w20181 = w20228 ^ w20189;
	assign w20188 = w20218 ^ w20181;
	assign w20264 = w20185 ^ w20188;
	assign w20260 = w20181 ^ w20182;
	assign w20258 = w20268 & w20297;
	assign w20252 = w20260 & w20293;
	assign w20237 = w20252 ^ w44219;
	assign w20213 = w20252 ^ w20255;
	assign w20210 = ~w20213;
	assign w20209 = w20252 ^ w20253;
	assign w20203 = w20248 ^ w20237;
	assign w20200 = ~w20203;
	assign w20197 = w20253 ^ w20237;
	assign w20251 = w20264 & w20296;
	assign w20229 = w20247 ^ w20251;
	assign w20207 = ~w20229;
	assign w20206 = w20207 ^ w20245;
	assign w20202 = w20206 ^ w44220;
	assign w20205 = w20244 ^ w20202;
	assign w20249 = w20268 & w20299;
	assign w20243 = w20260 & w20308;
	assign w20242 = w20264 & w20305;
	assign w20208 = w20253 ^ w20242;
	assign w20204 = ~w20208;
	assign w20309 = w20204 ^ w20205;
	assign w44218 = w20243 ^ w20244;
	assign w20225 = w20249 ^ w44218;
	assign w20226 = w20250 ^ w20225;
	assign w20230 = w20258 ^ w20226;
	assign w20235 = w20259 ^ w20230;
	assign w48906 = w44219 ^ w20235;
	assign w20310 = w20235 ^ w20209;
	assign w20201 = w20225 ^ w20202;
	assign w48904 = w20200 ^ w20201;
	assign w20199 = w20257 ^ w20230;
	assign w48905 = w20198 ^ w20199;
	assign w48907 = w20226 ^ w20197;
	assign w6952 = w48906 ^ w48905;
	assign w20212 = w20216 ^ w44218;
	assign w20215 = w44220 ^ w20212;
	assign w20312 = w20214 ^ w20215;
	assign w20211 = w20207 ^ w20212;
	assign w20311 = w20210 ^ w20211;
	assign w47572 = w48574 ^ w1914;
	assign w20431 = w47572 ^ w20432;
	assign w20358 = w47572 ^ w47566;
	assign w20428 = w20358 ^ w20353;
	assign w20435 = w20352 ^ w20358;
	assign w20433 = w20368 ^ w20435;
	assign w20438 = w47567 ^ w20358;
	assign w20434 = w47571 ^ w20438;
	assign w20437 = w47572 ^ w20313;
	assign w20424 = w20433 & w20431;
	assign w20375 = w20418 ^ w20424;
	assign w20416 = w20375 ^ w20366;
	assign w20423 = w47572 & w20437;
	assign w20421 = w20438 & w20434;
	assign w20415 = w20421 ^ w20373;
	assign w20420 = w20435 & w20428;
	assign w20412 = w20416 & w20415;
	assign w44222 = w20417 ^ w20420;
	assign w20330 = w20356 ^ w44222;
	assign w20414 = w20330 ^ w20355;
	assign w20411 = w20412 ^ w20414;
	assign w20370 = w20418 ^ w44222;
	assign w20326 = w20421 ^ w20370;
	assign w20408 = w47571 ^ w20326;
	assign w44225 = w20417 ^ w20423;
	assign w20329 = w20361 ^ w44225;
	assign w20372 = w47567 ^ w20329;
	assign w20407 = w20412 ^ w20372;
	assign w20406 = w20407 & w20408;
	assign w20405 = w20406 ^ w20414;
	assign w20404 = w20412 ^ w20406;
	assign w20325 = w20406 ^ w20370;
	assign w20324 = w20406 ^ w20423;
	assign w20319 = w20324 ^ w20420;
	assign w20403 = w20414 & w20404;
	assign w20401 = w20403 ^ w20411;
	assign w20391 = w20405 & w47572;
	assign w20382 = w20405 & w20437;
	assign w44224 = w20403 ^ w20421;
	assign w20395 = w44224 ^ w20373;
	assign w20393 = w20395 & w20432;
	assign w20384 = w20395 & w20436;
	assign w20362 = w47571 ^ w44224;
	assign w20402 = w20362 ^ w20325;
	assign w20392 = w20402 & w20431;
	assign w20383 = w20402 & w20433;
	assign w20367 = w44225 ^ w20352;
	assign w20413 = w20375 ^ w20367;
	assign w20410 = w20413 & w20411;
	assign w20409 = w20410 ^ w20372;
	assign w20321 = w20410 ^ w20422;
	assign w20317 = w20321 ^ w20357;
	assign w20320 = w47565 ^ w20317;
	assign w20397 = w20319 ^ w20320;
	assign w20318 = w20410 ^ w20366;
	assign w20316 = w47567 ^ w20317;
	assign w20400 = w20409 & w20401;
	assign w20365 = w20400 ^ w20375;
	assign w20399 = w20365 ^ w20367;
	assign w20323 = w20400 ^ w20424;
	assign w20315 = w20362 ^ w20323;
	assign w20322 = w20352 ^ w20315;
	assign w20398 = w20319 ^ w20322;
	assign w20396 = w20365 ^ w20318;
	assign w20394 = w20315 ^ w20316;
	assign w20390 = w20396 & w20426;
	assign w20389 = w20399 & w20438;
	assign w20388 = w20409 & w20428;
	assign w20332 = w20388 ^ w20389;
	assign w20387 = w20397 & w20429;
	assign w20386 = w20394 & w20427;
	assign w20347 = w20386 ^ w20389;
	assign w20344 = ~w20347;
	assign w20343 = w20386 ^ w20387;
	assign w20385 = w20398 & w20430;
	assign w20381 = w20396 & w20441;
	assign w20363 = w20381 ^ w20385;
	assign w20348 = w20390 ^ w20381;
	assign w20341 = ~w20363;
	assign w20380 = w20399 & w20434;
	assign w20350 = w20388 ^ w20380;
	assign w20379 = w20409 & w20435;
	assign w20340 = w20341 ^ w20379;
	assign w20378 = w20397 & w20440;
	assign w20377 = w20394 & w20442;
	assign w20376 = w20398 & w20439;
	assign w20342 = w20387 ^ w20376;
	assign w20338 = ~w20342;
	assign w44223 = w20377 ^ w20378;
	assign w20359 = w20383 ^ w44223;
	assign w20360 = w20384 ^ w20359;
	assign w20364 = w20392 ^ w20360;
	assign w20369 = w20393 ^ w20364;
	assign w20444 = w20369 ^ w20343;
	assign w20333 = w20391 ^ w20364;
	assign w48860 = w20332 ^ w20333;
	assign w6909 = w48866 ^ w48860;
	assign w7180 = w48860 ^ w48865;
	assign w7044 = ~w7180;
	assign w20346 = w20350 ^ w44223;
	assign w20345 = w20341 ^ w20346;
	assign w20445 = w20344 ^ w20345;
	assign w44226 = w20389 ^ w20390;
	assign w48861 = w44226 ^ w20369;
	assign w7060 = w45271 ^ w48861;
	assign w20371 = w20386 ^ w44226;
	assign w20337 = w20382 ^ w20371;
	assign w20334 = ~w20337;
	assign w20331 = w20387 ^ w20371;
	assign w48862 = w20360 ^ w20331;
	assign w7148 = w48862 ^ w48867;
	assign w44227 = w20391 ^ w20393;
	assign w20349 = w44227 ^ w20346;
	assign w20446 = w20348 ^ w20349;
	assign w20336 = w20340 ^ w44227;
	assign w20339 = w20378 ^ w20336;
	assign w20443 = w20338 ^ w20339;
	assign w20335 = w20359 ^ w20336;
	assign w48859 = w20334 ^ w20335;
	assign w6906 = w6907 ^ w48859;
	assign w7183 = w48859 ^ w48864;
	assign w7036 = ~w7183;
	assign w44805 = w34353 ^ w34359;
	assign w34265 = w34297 ^ w44805;
	assign w34308 = w47559 ^ w34265;
	assign w34343 = w34348 ^ w34308;
	assign w34303 = w44805 ^ w34288;
	assign w34349 = w34311 ^ w34303;
	assign w44806 = w34353 ^ w34356;
	assign w34306 = w34354 ^ w44806;
	assign w34262 = w34357 ^ w34306;
	assign w34344 = w47563 ^ w34262;
	assign w34342 = w34343 & w34344;
	assign w34260 = w34342 ^ w34359;
	assign w34255 = w34260 ^ w34356;
	assign w34340 = w34348 ^ w34342;
	assign w34261 = w34342 ^ w34306;
	assign w34266 = w34292 ^ w44806;
	assign w34350 = w34266 ^ w34291;
	assign w34341 = w34342 ^ w34350;
	assign w34347 = w34348 ^ w34350;
	assign w34346 = w34349 & w34347;
	assign w34345 = w34346 ^ w34308;
	assign w34257 = w34346 ^ w34358;
	assign w34253 = w34257 ^ w34293;
	assign w34256 = w47557 ^ w34253;
	assign w34333 = w34255 ^ w34256;
	assign w34254 = w34346 ^ w34302;
	assign w34252 = w47559 ^ w34253;
	assign w34339 = w34350 & w34340;
	assign w34337 = w34339 ^ w34347;
	assign w34336 = w34345 & w34337;
	assign w34301 = w34336 ^ w34311;
	assign w34335 = w34301 ^ w34303;
	assign w34259 = w34336 ^ w34360;
	assign w34332 = w34301 ^ w34254;
	assign w34327 = w34341 & w47564;
	assign w34326 = w34332 & w34362;
	assign w34325 = w34335 & w34374;
	assign w34324 = w34345 & w34364;
	assign w34268 = w34324 ^ w34325;
	assign w34323 = w34333 & w34365;
	assign w34318 = w34341 & w34373;
	assign w34317 = w34332 & w34377;
	assign w34284 = w34326 ^ w34317;
	assign w34316 = w34335 & w34370;
	assign w34286 = w34324 ^ w34316;
	assign w34315 = w34345 & w34371;
	assign w34314 = w34333 & w34376;
	assign w44808 = w34325 ^ w34326;
	assign w44810 = w34339 ^ w34357;
	assign w34331 = w44810 ^ w34309;
	assign w34329 = w34331 & w34368;
	assign w44809 = w34327 ^ w34329;
	assign w34320 = w34331 & w34372;
	assign w34298 = w47563 ^ w44810;
	assign w34338 = w34298 ^ w34261;
	assign w34251 = w34298 ^ w34259;
	assign w34258 = w34288 ^ w34251;
	assign w34334 = w34255 ^ w34258;
	assign w34330 = w34251 ^ w34252;
	assign w34328 = w34338 & w34367;
	assign w34322 = w34330 & w34363;
	assign w34307 = w34322 ^ w44808;
	assign w34283 = w34322 ^ w34325;
	assign w34280 = ~w34283;
	assign w34279 = w34322 ^ w34323;
	assign w34273 = w34318 ^ w34307;
	assign w34270 = ~w34273;
	assign w34267 = w34323 ^ w34307;
	assign w34321 = w34334 & w34366;
	assign w34299 = w34317 ^ w34321;
	assign w34277 = ~w34299;
	assign w34276 = w34277 ^ w34315;
	assign w34272 = w34276 ^ w44809;
	assign w34275 = w34314 ^ w34272;
	assign w34319 = w34338 & w34369;
	assign w34313 = w34330 & w34378;
	assign w34312 = w34334 & w34375;
	assign w34278 = w34323 ^ w34312;
	assign w34274 = ~w34278;
	assign w34379 = w34274 ^ w34275;
	assign w7078 = w45446 ^ w34379;
	assign w48846 = ~w34379;
	assign w44807 = w34313 ^ w34314;
	assign w34295 = w34319 ^ w44807;
	assign w34296 = w34320 ^ w34295;
	assign w48848 = w34296 ^ w34267;
	assign w34300 = w34328 ^ w34296;
	assign w34269 = w34327 ^ w34300;
	assign w48844 = w34268 ^ w34269;
	assign w34305 = w34329 ^ w34300;
	assign w48845 = w44808 ^ w34305;
	assign w34380 = w34305 ^ w34279;
	assign w48847 = ~w34380;
	assign w6938 = w48851 ^ w48844;
	assign w7080 = w48852 ^ w48845;
	assign w7152 = w48848 ^ w48853;
	assign w7086 = ~w7152;
	assign w7076 = w45447 ^ w34380;
	assign w34271 = w34295 ^ w34272;
	assign w48843 = w34270 ^ w34271;
	assign w7190 = w48843 ^ w48850;
	assign w7073 = ~w7190;
	assign w34282 = w34286 ^ w44807;
	assign w34285 = w44809 ^ w34282;
	assign w34382 = w34284 ^ w34285;
	assign w34281 = w34277 ^ w34282;
	assign w34381 = w34280 ^ w34281;
	assign w7176 = w48861 ^ w48866;
	assign w7018 = ~w7176;
	assign w45450 = ~w20309;
	assign w45451 = ~w20310;
	assign w7100 = w45451 ^ w45450;
	assign w45452 = ~w20311;
	assign w45453 = ~w20312;
	assign w45454 = ~w20443;
	assign w7172 = w45454 ^ w45271;
	assign w45455 = ~w20444;
	assign w7039 = w48862 ^ w45455;
	assign w45456 = ~w20445;
	assign w7062 = w48864 ^ w45456;
	assign w7187 = w45456 ^ w48863;
	assign w45457 = ~w20446;
	assign w6903 = w13745 ^ w45457;
	assign w7188 = w45457 ^ w45273;
	assign w45792 = ~w34381;
	assign w7090 = w7086 ^ w45792;
	assign w7192 = w45792 ^ w48849;
	assign w45793 = ~w34382;
	assign w7191 = w45793 ^ w45448;
	assign w45904 = ~w6033;
	assign w6045 = w45904 ^ w45805;
	assign w6047 = w6046 ^ w6045;
	assign w48414 = ~w6047;
	assign w6050 = w45904 ^ w48503;
	assign w48416 = w6051 ^ w6050;
	assign w6230 = w45904 ^ w48494;
	assign w5961 = w6230 ^ w6229;
	assign w48417 = w5961 ^ w6017;
	assign w47659 = w48414 ^ w105;
	assign w34504 = w47659 ^ w34508;
	assign w34438 = w47659 ^ w47658;
	assign w34503 = w34438 ^ w34505;
	assign w34511 = w47653 ^ w47659;
	assign w34491 = w34508 & w34504;
	assign w47656 = w48417 ^ w108;
	assign w34424 = w47656 ^ w47654;
	assign w34510 = w47656 ^ w47653;
	assign w34506 = w34510 ^ w34438;
	assign w34512 = w47658 ^ w47656;
	assign w34497 = w34422 ^ w34512;
	assign w34384 = w34424 ^ w34422;
	assign w34383 = w34424 ^ w47655;
	assign w34507 = w47660 ^ w34383;
	assign w34493 = w47660 & w34507;
	assign w34488 = w34512 & w34497;
	assign w47657 = w48416 ^ w107;
	assign w34421 = w47659 ^ w47657;
	assign w34423 = w47658 ^ w34421;
	assign w34499 = w47654 ^ w34423;
	assign w34496 = w47655 ^ w34423;
	assign w34498 = w34428 ^ w34423;
	assign w34502 = w34421 ^ w34510;
	assign w34501 = w47660 ^ w34502;
	assign w34398 = w47657 ^ w47658;
	assign w34500 = w34421 ^ w34384;
	assign w34495 = w34502 & w34506;
	assign w34427 = w34495 ^ w34424;
	assign w34494 = w34503 & w34501;
	assign w34445 = w34488 ^ w34494;
	assign w34492 = w34511 & w34496;
	assign w34426 = w34492 ^ w34422;
	assign w34490 = w34505 & w34498;
	assign w34489 = w34510 & w34499;
	assign w34425 = w34489 ^ w34423;
	assign w34431 = w34427 ^ w34425;
	assign w34436 = w47653 ^ w34431;
	assign w34486 = w34445 ^ w34436;
	assign w34397 = w34488 ^ w34489;
	assign w34444 = w34397 ^ w34398;
	assign w34443 = w34444 ^ w34426;
	assign w34485 = w34491 ^ w34443;
	assign w34487 = w34509 & w34500;
	assign w34482 = w34486 & w34485;
	assign w44811 = w34487 ^ w34490;
	assign w34400 = w34426 ^ w44811;
	assign w34484 = w34400 ^ w34425;
	assign w34481 = w34482 ^ w34484;
	assign w34440 = w34488 ^ w44811;
	assign w34396 = w34491 ^ w34440;
	assign w34478 = w47659 ^ w34396;
	assign w44814 = w34487 ^ w34493;
	assign w34399 = w34431 ^ w44814;
	assign w34442 = w47655 ^ w34399;
	assign w34477 = w34482 ^ w34442;
	assign w34476 = w34477 & w34478;
	assign w34474 = w34482 ^ w34476;
	assign w34395 = w34476 ^ w34440;
	assign w34394 = w34476 ^ w34493;
	assign w34389 = w34394 ^ w34490;
	assign w34473 = w34484 & w34474;
	assign w34471 = w34473 ^ w34481;
	assign w44813 = w34473 ^ w34491;
	assign w34465 = w44813 ^ w34443;
	assign w34454 = w34465 & w34506;
	assign w34463 = w34465 & w34502;
	assign w34432 = w47659 ^ w44813;
	assign w34472 = w34432 ^ w34395;
	assign w34462 = w34472 & w34501;
	assign w34453 = w34472 & w34503;
	assign w34475 = w34476 ^ w34484;
	assign w34461 = w34475 & w47660;
	assign w34452 = w34475 & w34507;
	assign w34437 = w44814 ^ w34422;
	assign w34483 = w34445 ^ w34437;
	assign w34480 = w34483 & w34481;
	assign w34479 = w34480 ^ w34442;
	assign w34391 = w34480 ^ w34492;
	assign w34387 = w34391 ^ w34427;
	assign w34390 = w47653 ^ w34387;
	assign w34467 = w34389 ^ w34390;
	assign w34388 = w34480 ^ w34436;
	assign w34386 = w47655 ^ w34387;
	assign w34470 = w34479 & w34471;
	assign w34435 = w34470 ^ w34445;
	assign w34469 = w34435 ^ w34437;
	assign w34393 = w34470 ^ w34494;
	assign w34385 = w34432 ^ w34393;
	assign w34392 = w34422 ^ w34385;
	assign w34468 = w34389 ^ w34392;
	assign w34466 = w34435 ^ w34388;
	assign w34464 = w34385 ^ w34386;
	assign w34460 = w34466 & w34496;
	assign w34459 = w34469 & w34508;
	assign w34458 = w34479 & w34498;
	assign w34402 = w34458 ^ w34459;
	assign w34457 = w34467 & w34499;
	assign w34456 = w34464 & w34497;
	assign w34417 = w34456 ^ w34459;
	assign w34414 = ~w34417;
	assign w34413 = w34456 ^ w34457;
	assign w34455 = w34468 & w34500;
	assign w34451 = w34466 & w34511;
	assign w34433 = w34451 ^ w34455;
	assign w34418 = w34460 ^ w34451;
	assign w34411 = ~w34433;
	assign w34450 = w34469 & w34504;
	assign w34420 = w34458 ^ w34450;
	assign w34449 = w34479 & w34505;
	assign w34410 = w34411 ^ w34449;
	assign w34448 = w34467 & w34510;
	assign w34447 = w34464 & w34512;
	assign w34446 = w34468 & w34509;
	assign w34412 = w34457 ^ w34446;
	assign w34408 = ~w34412;
	assign w44812 = w34447 ^ w34448;
	assign w34429 = w34453 ^ w44812;
	assign w34430 = w34454 ^ w34429;
	assign w34434 = w34462 ^ w34430;
	assign w34403 = w34461 ^ w34434;
	assign w48664 = w34402 ^ w34403;
	assign w6428 = ~w48664;
	assign w6427 = w6428 ^ w48658;
	assign w6756 = w6426 ^ w6427;
	assign w48545 = w6756 ^ w6694;
	assign w47601 = w48545 ^ w1949;
	assign w6440 = w48668 ^ w6428;
	assign w6701 = w48659 ^ w48664;
	assign w6565 = ~w6701;
	assign w6563 = w6565 ^ w6689;
	assign w6543 = w6701 ^ w6699;
	assign w48569 = w6543 ^ w6544;
	assign w47577 = w48569 ^ w1973;
	assign w34439 = w34463 ^ w34434;
	assign w34514 = w34439 ^ w34413;
	assign w34416 = w34420 ^ w44812;
	assign w34415 = w34411 ^ w34416;
	assign w34515 = w34414 ^ w34415;
	assign w6556 = w45752 ^ w34515;
	assign w48662 = ~w34515;
	assign w6708 = w45477 ^ w48662;
	assign w6568 = w6708 ^ w6699;
	assign w48552 = w48658 ^ w6568;
	assign w47594 = w48552 ^ w1956;
	assign w6546 = w6708 ^ w6706;
	assign w48567 = w6546 ^ w6547;
	assign w47579 = w48567 ^ w1971;
	assign w31875 = w47579 ^ w47577;
	assign w6424 = w34515 ^ w45470;
	assign w6757 = w6423 ^ w6424;
	assign w48543 = w6757 ^ w6702;
	assign w47603 = w48543 ^ w1947;
	assign w20485 = w47603 ^ w47601;
	assign w44815 = w34459 ^ w34460;
	assign w48665 = w44815 ^ w34439;
	assign w6697 = w48660 ^ w48665;
	assign w6539 = ~w6697;
	assign w6536 = w6539 ^ w6694;
	assign w48570 = w6536 ^ w6537;
	assign w47576 = w48570 ^ w1974;
	assign w6562 = w6697 ^ w6684;
	assign w48555 = w45475 ^ w6562;
	assign w47591 = w48555 ^ w1959;
	assign w6430 = w48665 ^ w48659;
	assign w6755 = w6429 ^ w6430;
	assign w48546 = w6755 ^ w6689;
	assign w47600 = w48546 ^ w1950;
	assign w6553 = w6538 ^ w48665;
	assign w34441 = w34456 ^ w44815;
	assign w34407 = w34452 ^ w34441;
	assign w34404 = ~w34407;
	assign w34401 = w34457 ^ w34441;
	assign w48666 = w34430 ^ w34401;
	assign w6669 = w48661 ^ w48666;
	assign w6676 = w48666 ^ w48670;
	assign w6532 = w6669 ^ w45567;
	assign w48573 = w6532 ^ w6533;
	assign w6572 = w6706 ^ w6669;
	assign w6441 = ~w6676;
	assign w48550 = w45470 ^ w6572;
	assign w47596 = w48550 ^ w1954;
	assign w6439 = w6441 ^ w48673;
	assign w6750 = w6439 ^ w6440;
	assign w48562 = w6750 ^ w6697;
	assign w6437 = w6676 ^ w48672;
	assign w6435 = w6676 ^ w45568;
	assign w47573 = w48573 ^ w1977;
	assign w31964 = w47576 ^ w47573;
	assign w31956 = w31875 ^ w31964;
	assign w31965 = w47573 ^ w47579;
	assign w47584 = w48562 ^ w1966;
	assign w44816 = w34461 ^ w34463;
	assign w34419 = w44816 ^ w34416;
	assign w34516 = w34418 ^ w34419;
	assign w34406 = w34410 ^ w44816;
	assign w34409 = w34448 ^ w34406;
	assign w34513 = w34408 ^ w34409;
	assign w34405 = w34429 ^ w34406;
	assign w48663 = w34404 ^ w34405;
	assign w6438 = w48667 ^ w48663;
	assign w6583 = w48663 ^ w45477;
	assign w6751 = w6437 ^ w6438;
	assign w48561 = w6751 ^ w6701;
	assign w47585 = w48561 ^ w1965;
	assign w48544 = w6582 ^ w6583;
	assign w47602 = w48544 ^ w1948;
	assign w20487 = w47602 ^ w20485;
	assign w20502 = w47603 ^ w47602;
	assign w20576 = w47602 ^ w47600;
	assign w20462 = w47601 ^ w47602;
	assign w6704 = w48658 ^ w48663;
	assign w6557 = ~w6704;
	assign w6545 = w6704 ^ w6702;
	assign w6566 = w6557 ^ w6694;
	assign w48568 = w48667 ^ w6545;
	assign w47578 = w48568 ^ w1972;
	assign w31877 = w47578 ^ w31875;
	assign w31892 = w47579 ^ w47578;
	assign w31960 = w31964 ^ w31892;
	assign w31966 = w47578 ^ w47576;
	assign w31852 = w47577 ^ w47578;
	assign w31963 = w47573 ^ w47578;
	assign w31949 = w31956 & w31960;
	assign w48549 = w48666 ^ w6577;
	assign w47597 = w48549 ^ w1953;
	assign w20574 = w47600 ^ w47597;
	assign w20570 = w20574 ^ w20502;
	assign w20566 = w20485 ^ w20574;
	assign w20575 = w47597 ^ w47603;
	assign w20573 = w47597 ^ w47602;
	assign w20559 = w20566 & w20570;
	assign w6555 = w6557 ^ w48671;
	assign w48560 = w6555 ^ w6556;
	assign w47586 = w48560 ^ w1964;
	assign w25400 = w47586 ^ w47584;
	assign w25286 = w47585 ^ w47586;
	assign w45790 = ~w34514;
	assign w6686 = w45790 ^ w45751;
	assign w6578 = w6686 ^ w45567;
	assign w48548 = w6578 ^ w6579;
	assign w6549 = w6686 ^ w6669;
	assign w47598 = w48548 ^ w1952;
	assign w20563 = w47598 ^ w20487;
	assign w20488 = w47600 ^ w47598;
	assign w20491 = w20559 ^ w20488;
	assign w20553 = w20574 & w20563;
	assign w20489 = w20553 ^ w20487;
	assign w20495 = w20491 ^ w20489;
	assign w20500 = w47597 ^ w20495;
	assign w6534 = w6686 ^ w6684;
	assign w48572 = w45476 ^ w6534;
	assign w47574 = w48572 ^ w1976;
	assign w31953 = w47574 ^ w31877;
	assign w31878 = w47576 ^ w47574;
	assign w31881 = w31949 ^ w31878;
	assign w31943 = w31964 & w31953;
	assign w31879 = w31943 ^ w31877;
	assign w31885 = w31881 ^ w31879;
	assign w31890 = w47573 ^ w31885;
	assign w48565 = w48674 ^ w6549;
	assign w47581 = w48565 ^ w1969;
	assign w25398 = w47584 ^ w47581;
	assign w25397 = w47581 ^ w47586;
	assign w6559 = w6668 ^ w45790;
	assign w48557 = w6559 ^ w6560;
	assign w47589 = w48557 ^ w1961;
	assign w13786 = w47591 ^ w47589;
	assign w13873 = w47589 ^ w47594;
	assign w45791 = ~w34516;
	assign w48542 = w45791 ^ w6584;
	assign w47604 = w48542 ^ w1946;
	assign w20565 = w47604 ^ w20566;
	assign w20492 = w47604 ^ w47598;
	assign w20562 = w20492 ^ w20487;
	assign w6709 = w45470 ^ w45791;
	assign w6548 = w6709 ^ w6668;
	assign w48566 = w45753 ^ w6548;
	assign w47580 = w48566 ^ w1970;
	assign w31955 = w47580 ^ w31956;
	assign w31882 = w47580 ^ w47574;
	assign w31952 = w31882 ^ w31877;
	assign w6436 = w45753 ^ w45791;
	assign w6570 = w6709 ^ w6702;
	assign w6558 = w6709 ^ w6676;
	assign w48558 = w45569 ^ w6558;
	assign w47588 = w48558 ^ w1962;
	assign w6752 = w6435 ^ w6436;
	assign w48559 = w6752 ^ w6708;
	assign w47587 = w48559 ^ w1963;
	assign w25309 = w47587 ^ w47585;
	assign w25311 = w47586 ^ w25309;
	assign w25390 = w25309 ^ w25398;
	assign w25389 = w47588 ^ w25390;
	assign w25326 = w47587 ^ w47586;
	assign w25394 = w25398 ^ w25326;
	assign w25399 = w47581 ^ w47587;
	assign w25383 = w25390 & w25394;
	assign w45797 = ~w34513;
	assign w6581 = w45797 ^ w48660;
	assign w48547 = w6580 ^ w6581;
	assign w6551 = w45790 ^ w45797;
	assign w48564 = w6550 ^ w6551;
	assign w47599 = w48547 ^ w1951;
	assign w20560 = w47599 ^ w20487;
	assign w20486 = w47599 ^ w47597;
	assign w20561 = w20486 ^ w20576;
	assign w20569 = w20486 ^ w20492;
	assign w20567 = w20502 ^ w20569;
	assign w20572 = w47599 ^ w20492;
	assign w20568 = w47603 ^ w20572;
	assign w20448 = w20488 ^ w20486;
	assign w20564 = w20485 ^ w20448;
	assign w20447 = w20488 ^ w47599;
	assign w20571 = w47604 ^ w20447;
	assign w20558 = w20567 & w20565;
	assign w20557 = w47604 & w20571;
	assign w20556 = w20575 & w20560;
	assign w20490 = w20556 ^ w20486;
	assign w20555 = w20572 & w20568;
	assign w20554 = w20569 & w20562;
	assign w20552 = w20576 & w20561;
	assign w20509 = w20552 ^ w20558;
	assign w20550 = w20509 ^ w20500;
	assign w20461 = w20552 ^ w20553;
	assign w20508 = w20461 ^ w20462;
	assign w20507 = w20508 ^ w20490;
	assign w20549 = w20555 ^ w20507;
	assign w20551 = w20573 & w20564;
	assign w20546 = w20550 & w20549;
	assign w6693 = w45475 ^ w45797;
	assign w6554 = w6693 ^ w45566;
	assign w6535 = w6693 ^ w6689;
	assign w6552 = ~w6554;
	assign w48563 = w6552 ^ w6553;
	assign w47583 = w48563 ^ w1967;
	assign w25384 = w47583 ^ w25311;
	assign w25310 = w47583 ^ w47581;
	assign w25385 = w25310 ^ w25400;
	assign w25380 = w25399 & w25384;
	assign w25314 = w25380 ^ w25310;
	assign w25376 = w25400 & w25385;
	assign w48571 = w45750 ^ w6535;
	assign w47575 = w48571 ^ w1975;
	assign w31950 = w47575 ^ w31877;
	assign w31876 = w47575 ^ w47573;
	assign w31951 = w31876 ^ w31966;
	assign w31959 = w31876 ^ w31882;
	assign w31957 = w31892 ^ w31959;
	assign w31962 = w47575 ^ w31882;
	assign w31958 = w47579 ^ w31962;
	assign w31838 = w31878 ^ w31876;
	assign w31954 = w31875 ^ w31838;
	assign w31837 = w31878 ^ w47575;
	assign w31961 = w47580 ^ w31837;
	assign w31948 = w31957 & w31955;
	assign w31947 = w47580 & w31961;
	assign w31946 = w31965 & w31950;
	assign w31880 = w31946 ^ w31876;
	assign w31945 = w31962 & w31958;
	assign w31944 = w31959 & w31952;
	assign w31942 = w31966 & w31951;
	assign w31899 = w31942 ^ w31948;
	assign w31940 = w31899 ^ w31890;
	assign w31851 = w31942 ^ w31943;
	assign w31898 = w31851 ^ w31852;
	assign w31897 = w31898 ^ w31880;
	assign w31939 = w31945 ^ w31897;
	assign w31941 = w31963 & w31954;
	assign w31936 = w31940 & w31939;
	assign w6561 = w6693 ^ w6687;
	assign w47582 = w48564 ^ w1968;
	assign w25387 = w47582 ^ w25311;
	assign w25312 = w47584 ^ w47582;
	assign w25315 = w25383 ^ w25312;
	assign w25316 = w47588 ^ w47582;
	assign w25386 = w25316 ^ w25311;
	assign w25393 = w25310 ^ w25316;
	assign w25391 = w25326 ^ w25393;
	assign w25396 = w47583 ^ w25316;
	assign w25392 = w47587 ^ w25396;
	assign w25272 = w25312 ^ w25310;
	assign w25388 = w25309 ^ w25272;
	assign w25271 = w25312 ^ w47583;
	assign w25395 = w47588 ^ w25271;
	assign w25382 = w25391 & w25389;
	assign w25333 = w25376 ^ w25382;
	assign w25381 = w47588 & w25395;
	assign w25379 = w25396 & w25392;
	assign w25378 = w25393 & w25386;
	assign w25377 = w25398 & w25387;
	assign w25313 = w25377 ^ w25311;
	assign w25319 = w25315 ^ w25313;
	assign w25324 = w47581 ^ w25319;
	assign w25374 = w25333 ^ w25324;
	assign w25285 = w25376 ^ w25377;
	assign w25332 = w25285 ^ w25286;
	assign w25331 = w25332 ^ w25314;
	assign w25373 = w25379 ^ w25331;
	assign w25375 = w25397 & w25388;
	assign w25370 = w25374 & w25373;
	assign w48556 = w45751 ^ w6561;
	assign w47590 = w48556 ^ w1960;
	assign w13792 = w47596 ^ w47590;
	assign w13869 = w13786 ^ w13792;
	assign w13872 = w47591 ^ w13792;
	assign w44228 = w20551 ^ w20557;
	assign w20501 = w44228 ^ w20486;
	assign w20547 = w20509 ^ w20501;
	assign w20463 = w20495 ^ w44228;
	assign w20506 = w47599 ^ w20463;
	assign w20541 = w20546 ^ w20506;
	assign w44229 = w20551 ^ w20554;
	assign w20504 = w20552 ^ w44229;
	assign w20460 = w20555 ^ w20504;
	assign w20542 = w47603 ^ w20460;
	assign w20540 = w20541 & w20542;
	assign w20538 = w20546 ^ w20540;
	assign w20459 = w20540 ^ w20504;
	assign w20458 = w20540 ^ w20557;
	assign w20453 = w20458 ^ w20554;
	assign w20464 = w20490 ^ w44229;
	assign w20548 = w20464 ^ w20489;
	assign w20539 = w20540 ^ w20548;
	assign w20545 = w20546 ^ w20548;
	assign w20544 = w20547 & w20545;
	assign w20543 = w20544 ^ w20506;
	assign w20455 = w20544 ^ w20556;
	assign w20451 = w20455 ^ w20491;
	assign w20454 = w47597 ^ w20451;
	assign w20531 = w20453 ^ w20454;
	assign w20452 = w20544 ^ w20500;
	assign w20450 = w47599 ^ w20451;
	assign w20537 = w20548 & w20538;
	assign w20535 = w20537 ^ w20545;
	assign w20534 = w20543 & w20535;
	assign w20499 = w20534 ^ w20509;
	assign w20533 = w20499 ^ w20501;
	assign w20457 = w20534 ^ w20558;
	assign w20530 = w20499 ^ w20452;
	assign w20525 = w20539 & w47604;
	assign w20524 = w20530 & w20560;
	assign w20523 = w20533 & w20572;
	assign w20522 = w20543 & w20562;
	assign w20466 = w20522 ^ w20523;
	assign w20521 = w20531 & w20563;
	assign w20516 = w20539 & w20571;
	assign w20515 = w20530 & w20575;
	assign w20482 = w20524 ^ w20515;
	assign w20514 = w20533 & w20568;
	assign w20484 = w20522 ^ w20514;
	assign w20513 = w20543 & w20569;
	assign w20512 = w20531 & w20574;
	assign w44230 = w20523 ^ w20524;
	assign w44232 = w20537 ^ w20555;
	assign w20496 = w47603 ^ w44232;
	assign w20449 = w20496 ^ w20457;
	assign w20456 = w20486 ^ w20449;
	assign w20532 = w20453 ^ w20456;
	assign w20528 = w20449 ^ w20450;
	assign w20520 = w20528 & w20561;
	assign w20505 = w20520 ^ w44230;
	assign w20481 = w20520 ^ w20523;
	assign w20478 = ~w20481;
	assign w20477 = w20520 ^ w20521;
	assign w20465 = w20521 ^ w20505;
	assign w20519 = w20532 & w20564;
	assign w20471 = w20516 ^ w20505;
	assign w20468 = ~w20471;
	assign w20497 = w20515 ^ w20519;
	assign w20475 = ~w20497;
	assign w20474 = w20475 ^ w20513;
	assign w20536 = w20496 ^ w20459;
	assign w20517 = w20536 & w20567;
	assign w20526 = w20536 & w20565;
	assign w20511 = w20528 & w20576;
	assign w20510 = w20532 & w20573;
	assign w20476 = w20521 ^ w20510;
	assign w20472 = ~w20476;
	assign w43555 = w20511 ^ w20512;
	assign w20493 = w20517 ^ w43555;
	assign w20480 = w20484 ^ w43555;
	assign w20479 = w20475 ^ w20480;
	assign w20579 = w20478 ^ w20479;
	assign w20529 = w44232 ^ w20507;
	assign w20527 = w20529 & w20566;
	assign w20518 = w20529 & w20570;
	assign w20494 = w20518 ^ w20493;
	assign w20498 = w20526 ^ w20494;
	assign w20503 = w20527 ^ w20498;
	assign w48841 = w44230 ^ w20503;
	assign w20578 = w20503 ^ w20477;
	assign w20467 = w20525 ^ w20498;
	assign w48840 = w20466 ^ w20467;
	assign w48842 = w20494 ^ w20465;
	assign w7151 = w48842 ^ w48848;
	assign w6941 = w7151 ^ w48840;
	assign w7206 = w48841 ^ w48845;
	assign w7215 = w48840 ^ w48844;
	assign w7084 = w7215 ^ w7073;
	assign w7097 = ~w7215;
	assign w44231 = w20525 ^ w20527;
	assign w20483 = w44231 ^ w20480;
	assign w20580 = w20482 ^ w20483;
	assign w20470 = w20474 ^ w44231;
	assign w20473 = w20512 ^ w20470;
	assign w20577 = w20472 ^ w20473;
	assign w20469 = w20493 ^ w20470;
	assign w48839 = w20468 ^ w20469;
	assign w6942 = w48839 ^ w48843;
	assign w7220 = w6941 ^ w6942;
	assign w7071 = w7073 ^ w48839;
	assign w44430 = w25375 ^ w25381;
	assign w25325 = w44430 ^ w25310;
	assign w25371 = w25333 ^ w25325;
	assign w25287 = w25319 ^ w44430;
	assign w25330 = w47583 ^ w25287;
	assign w25365 = w25370 ^ w25330;
	assign w44431 = w25375 ^ w25378;
	assign w25328 = w25376 ^ w44431;
	assign w25284 = w25379 ^ w25328;
	assign w25366 = w47587 ^ w25284;
	assign w25364 = w25365 & w25366;
	assign w25362 = w25370 ^ w25364;
	assign w25283 = w25364 ^ w25328;
	assign w25282 = w25364 ^ w25381;
	assign w25277 = w25282 ^ w25378;
	assign w25288 = w25314 ^ w44431;
	assign w25372 = w25288 ^ w25313;
	assign w25363 = w25364 ^ w25372;
	assign w25369 = w25370 ^ w25372;
	assign w25368 = w25371 & w25369;
	assign w25367 = w25368 ^ w25330;
	assign w25279 = w25368 ^ w25380;
	assign w25275 = w25279 ^ w25315;
	assign w25278 = w47581 ^ w25275;
	assign w25355 = w25277 ^ w25278;
	assign w25276 = w25368 ^ w25324;
	assign w25274 = w47583 ^ w25275;
	assign w25361 = w25372 & w25362;
	assign w25359 = w25361 ^ w25369;
	assign w25358 = w25367 & w25359;
	assign w25323 = w25358 ^ w25333;
	assign w25357 = w25323 ^ w25325;
	assign w25281 = w25358 ^ w25382;
	assign w25354 = w25323 ^ w25276;
	assign w25349 = w25363 & w47588;
	assign w25348 = w25354 & w25384;
	assign w25347 = w25357 & w25396;
	assign w25346 = w25367 & w25386;
	assign w25290 = w25346 ^ w25347;
	assign w25345 = w25355 & w25387;
	assign w25340 = w25363 & w25395;
	assign w25339 = w25354 & w25399;
	assign w25306 = w25348 ^ w25339;
	assign w25338 = w25357 & w25392;
	assign w25308 = w25346 ^ w25338;
	assign w25337 = w25367 & w25393;
	assign w25336 = w25355 & w25398;
	assign w44432 = w25347 ^ w25348;
	assign w44434 = w25361 ^ w25379;
	assign w25320 = w47587 ^ w44434;
	assign w25360 = w25320 ^ w25283;
	assign w25350 = w25360 & w25389;
	assign w25341 = w25360 & w25391;
	assign w25273 = w25320 ^ w25281;
	assign w25352 = w25273 ^ w25274;
	assign w25344 = w25352 & w25385;
	assign w25329 = w25344 ^ w44432;
	assign w25305 = w25344 ^ w25347;
	assign w25302 = ~w25305;
	assign w25301 = w25344 ^ w25345;
	assign w25289 = w25345 ^ w25329;
	assign w25295 = w25340 ^ w25329;
	assign w25292 = ~w25295;
	assign w25335 = w25352 & w25400;
	assign w43569 = w25335 ^ w25336;
	assign w25304 = w25308 ^ w43569;
	assign w25317 = w25341 ^ w43569;
	assign w25280 = w25310 ^ w25273;
	assign w25356 = w25277 ^ w25280;
	assign w25334 = w25356 & w25397;
	assign w25300 = w25345 ^ w25334;
	assign w25296 = ~w25300;
	assign w25343 = w25356 & w25388;
	assign w25321 = w25339 ^ w25343;
	assign w25299 = ~w25321;
	assign w25298 = w25299 ^ w25337;
	assign w25303 = w25299 ^ w25304;
	assign w25403 = w25302 ^ w25303;
	assign w25353 = w44434 ^ w25331;
	assign w25351 = w25353 & w25390;
	assign w25342 = w25353 & w25394;
	assign w25318 = w25342 ^ w25317;
	assign w25322 = w25350 ^ w25318;
	assign w25327 = w25351 ^ w25322;
	assign w48889 = w44432 ^ w25327;
	assign w25402 = w25327 ^ w25301;
	assign w25291 = w25349 ^ w25322;
	assign w48888 = w25290 ^ w25291;
	assign w48890 = w25318 ^ w25289;
	assign w44433 = w25349 ^ w25351;
	assign w25307 = w44433 ^ w25304;
	assign w25404 = w25306 ^ w25307;
	assign w25294 = w25298 ^ w44433;
	assign w25297 = w25336 ^ w25294;
	assign w25401 = w25296 ^ w25297;
	assign w25293 = w25317 ^ w25294;
	assign w48887 = w25292 ^ w25293;
	assign w44705 = w31941 ^ w31947;
	assign w31853 = w31885 ^ w44705;
	assign w31896 = w47575 ^ w31853;
	assign w31931 = w31936 ^ w31896;
	assign w31891 = w44705 ^ w31876;
	assign w31937 = w31899 ^ w31891;
	assign w44706 = w31941 ^ w31944;
	assign w31894 = w31942 ^ w44706;
	assign w31850 = w31945 ^ w31894;
	assign w31932 = w47579 ^ w31850;
	assign w31930 = w31931 & w31932;
	assign w31848 = w31930 ^ w31947;
	assign w31843 = w31848 ^ w31944;
	assign w31928 = w31936 ^ w31930;
	assign w31849 = w31930 ^ w31894;
	assign w31854 = w31880 ^ w44706;
	assign w31938 = w31854 ^ w31879;
	assign w31929 = w31930 ^ w31938;
	assign w31935 = w31936 ^ w31938;
	assign w31934 = w31937 & w31935;
	assign w31933 = w31934 ^ w31896;
	assign w31845 = w31934 ^ w31946;
	assign w31841 = w31845 ^ w31881;
	assign w31844 = w47573 ^ w31841;
	assign w31921 = w31843 ^ w31844;
	assign w31842 = w31934 ^ w31890;
	assign w31840 = w47575 ^ w31841;
	assign w31927 = w31938 & w31928;
	assign w31925 = w31927 ^ w31935;
	assign w31924 = w31933 & w31925;
	assign w31889 = w31924 ^ w31899;
	assign w31923 = w31889 ^ w31891;
	assign w31847 = w31924 ^ w31948;
	assign w31920 = w31889 ^ w31842;
	assign w31915 = w31929 & w47580;
	assign w31914 = w31920 & w31950;
	assign w31913 = w31923 & w31962;
	assign w31912 = w31933 & w31952;
	assign w31856 = w31912 ^ w31913;
	assign w31911 = w31921 & w31953;
	assign w31906 = w31929 & w31961;
	assign w31905 = w31920 & w31965;
	assign w31872 = w31914 ^ w31905;
	assign w31904 = w31923 & w31958;
	assign w31874 = w31912 ^ w31904;
	assign w31903 = w31933 & w31959;
	assign w31902 = w31921 & w31964;
	assign w44708 = w31913 ^ w31914;
	assign w44710 = w31927 ^ w31945;
	assign w31919 = w44710 ^ w31897;
	assign w31917 = w31919 & w31956;
	assign w44709 = w31915 ^ w31917;
	assign w31908 = w31919 & w31960;
	assign w31886 = w47579 ^ w44710;
	assign w31926 = w31886 ^ w31849;
	assign w31839 = w31886 ^ w31847;
	assign w31846 = w31876 ^ w31839;
	assign w31922 = w31843 ^ w31846;
	assign w31918 = w31839 ^ w31840;
	assign w31916 = w31926 & w31955;
	assign w31910 = w31918 & w31951;
	assign w31895 = w31910 ^ w44708;
	assign w31871 = w31910 ^ w31913;
	assign w31868 = ~w31871;
	assign w31867 = w31910 ^ w31911;
	assign w31861 = w31906 ^ w31895;
	assign w31858 = ~w31861;
	assign w31855 = w31911 ^ w31895;
	assign w31909 = w31922 & w31954;
	assign w31887 = w31905 ^ w31909;
	assign w31865 = ~w31887;
	assign w31864 = w31865 ^ w31903;
	assign w31860 = w31864 ^ w44709;
	assign w31863 = w31902 ^ w31860;
	assign w31907 = w31926 & w31957;
	assign w31901 = w31918 & w31966;
	assign w31900 = w31922 & w31963;
	assign w31866 = w31911 ^ w31900;
	assign w31862 = ~w31866;
	assign w31967 = w31862 ^ w31863;
	assign w44707 = w31901 ^ w31902;
	assign w31883 = w31907 ^ w44707;
	assign w31859 = w31883 ^ w31860;
	assign w48872 = w31858 ^ w31859;
	assign w7034 = w7036 ^ w48872;
	assign w31884 = w31908 ^ w31883;
	assign w48875 = w31884 ^ w31855;
	assign w31888 = w31916 ^ w31884;
	assign w31857 = w31915 ^ w31888;
	assign w48873 = w31856 ^ w31857;
	assign w31893 = w31917 ^ w31888;
	assign w31968 = w31893 ^ w31867;
	assign w7157 = w48862 ^ w48875;
	assign w6908 = w7157 ^ w48873;
	assign w7234 = w6908 ^ w6909;
	assign w6904 = ~w7157;
	assign w6905 = w6904 ^ w48872;
	assign w7235 = w6905 ^ w6906;
	assign w48874 = w44708 ^ w31893;
	assign w31870 = w31874 ^ w44707;
	assign w31873 = w44709 ^ w31870;
	assign w31970 = w31872 ^ w31873;
	assign w31869 = w31865 ^ w31870;
	assign w31969 = w31868 ^ w31869;
	assign w45458 = ~w20577;
	assign w7203 = w45458 ^ w48846;
	assign w45459 = ~w20578;
	assign w7201 = w45459 ^ w48847;
	assign w45460 = ~w20579;
	assign w6944 = w45460 ^ w45448;
	assign w7125 = w45460 ^ w6947;
	assign w45461 = ~w20580;
	assign w6940 = w20177 ^ w45461;
	assign w45554 = ~w25402;
	assign w45555 = ~w25403;
	assign w45556 = ~w25404;
	assign w45561 = ~w25401;
	assign w45738 = ~w31967;
	assign w7033 = w7172 ^ w45738;
	assign w7031 = ~w7033;
	assign w7058 = w45738 ^ w45454;
	assign w45739 = ~w31968;
	assign w7011 = w7148 ^ w45739;
	assign w7166 = w45455 ^ w45739;
	assign w7040 = w7172 ^ w7166;
	assign w45740 = ~w31969;
	assign w45741 = ~w31970;
	assign w6902 = w6904 ^ w45741;
	assign w7236 = w6902 ^ w6903;
	assign w45905 = ~w6667;
	assign w6484 = w45905 ^ w48687;
	assign w6489 = w45905 ^ w45481;
	assign w48599 = w6488 ^ w6489;
	assign w6481 = w45905 ^ w48688;
	assign w48602 = w6480 ^ w6481;
	assign w47544 = w48602 ^ w1942;
	assign w31744 = w47544 ^ w47542;
	assign w31830 = w47544 ^ w47541;
	assign w31832 = w47546 ^ w47544;
	assign w31817 = w31742 ^ w31832;
	assign w31704 = w31744 ^ w31742;
	assign w31703 = w31744 ^ w47543;
	assign w31827 = w47548 ^ w31703;
	assign w31813 = w47548 & w31827;
	assign w31808 = w31832 & w31817;
	assign w48601 = w6483 ^ w6484;
	assign w47545 = w48601 ^ w1941;
	assign w31718 = w47545 ^ w47546;
	assign w47547 = w48599 ^ w1939;
	assign w31741 = w47547 ^ w47545;
	assign w31743 = w47546 ^ w31741;
	assign w31819 = w47542 ^ w31743;
	assign w31816 = w47543 ^ w31743;
	assign w31818 = w31748 ^ w31743;
	assign w31824 = w47547 ^ w31828;
	assign w31822 = w31741 ^ w31830;
	assign w31821 = w47548 ^ w31822;
	assign w31758 = w47547 ^ w47546;
	assign w31823 = w31758 ^ w31825;
	assign w31826 = w31830 ^ w31758;
	assign w31820 = w31741 ^ w31704;
	assign w31831 = w47541 ^ w47547;
	assign w31815 = w31822 & w31826;
	assign w31747 = w31815 ^ w31744;
	assign w31814 = w31823 & w31821;
	assign w31765 = w31808 ^ w31814;
	assign w31812 = w31831 & w31816;
	assign w31746 = w31812 ^ w31742;
	assign w31811 = w31828 & w31824;
	assign w31810 = w31825 & w31818;
	assign w31809 = w31830 & w31819;
	assign w31745 = w31809 ^ w31743;
	assign w31751 = w31747 ^ w31745;
	assign w31756 = w47541 ^ w31751;
	assign w31806 = w31765 ^ w31756;
	assign w31717 = w31808 ^ w31809;
	assign w31764 = w31717 ^ w31718;
	assign w31763 = w31764 ^ w31746;
	assign w31805 = w31811 ^ w31763;
	assign w31807 = w31829 & w31820;
	assign w31802 = w31806 & w31805;
	assign w44700 = w31807 ^ w31813;
	assign w31757 = w44700 ^ w31742;
	assign w31803 = w31765 ^ w31757;
	assign w31719 = w31751 ^ w44700;
	assign w31762 = w47543 ^ w31719;
	assign w31797 = w31802 ^ w31762;
	assign w44701 = w31807 ^ w31810;
	assign w31760 = w31808 ^ w44701;
	assign w31716 = w31811 ^ w31760;
	assign w31798 = w47547 ^ w31716;
	assign w31796 = w31797 & w31798;
	assign w31715 = w31796 ^ w31760;
	assign w31714 = w31796 ^ w31813;
	assign w31709 = w31714 ^ w31810;
	assign w31794 = w31802 ^ w31796;
	assign w31720 = w31746 ^ w44701;
	assign w31804 = w31720 ^ w31745;
	assign w31795 = w31796 ^ w31804;
	assign w31801 = w31802 ^ w31804;
	assign w31800 = w31803 & w31801;
	assign w31799 = w31800 ^ w31762;
	assign w31711 = w31800 ^ w31812;
	assign w31707 = w31711 ^ w31747;
	assign w31710 = w47541 ^ w31707;
	assign w31787 = w31709 ^ w31710;
	assign w31708 = w31800 ^ w31756;
	assign w31706 = w47543 ^ w31707;
	assign w31793 = w31804 & w31794;
	assign w31791 = w31793 ^ w31801;
	assign w31790 = w31799 & w31791;
	assign w31755 = w31790 ^ w31765;
	assign w31789 = w31755 ^ w31757;
	assign w31713 = w31790 ^ w31814;
	assign w31786 = w31755 ^ w31708;
	assign w31781 = w31795 & w47548;
	assign w31780 = w31786 & w31816;
	assign w31779 = w31789 & w31828;
	assign w31778 = w31799 & w31818;
	assign w31722 = w31778 ^ w31779;
	assign w31777 = w31787 & w31819;
	assign w31772 = w31795 & w31827;
	assign w31771 = w31786 & w31831;
	assign w31738 = w31780 ^ w31771;
	assign w31770 = w31789 & w31824;
	assign w31740 = w31778 ^ w31770;
	assign w31769 = w31799 & w31825;
	assign w31768 = w31787 & w31830;
	assign w44702 = w31779 ^ w31780;
	assign w44704 = w31793 ^ w31811;
	assign w31752 = w47547 ^ w44704;
	assign w31792 = w31752 ^ w31715;
	assign w31773 = w31792 & w31823;
	assign w31782 = w31792 & w31821;
	assign w31705 = w31752 ^ w31713;
	assign w31712 = w31742 ^ w31705;
	assign w31788 = w31709 ^ w31712;
	assign w31775 = w31788 & w31820;
	assign w31753 = w31771 ^ w31775;
	assign w31731 = ~w31753;
	assign w31730 = w31731 ^ w31769;
	assign w31784 = w31705 ^ w31706;
	assign w31767 = w31784 & w31832;
	assign w31766 = w31788 & w31829;
	assign w31732 = w31777 ^ w31766;
	assign w31728 = ~w31732;
	assign w43587 = w31767 ^ w31768;
	assign w31749 = w31773 ^ w43587;
	assign w31736 = w31740 ^ w43587;
	assign w31735 = w31731 ^ w31736;
	assign w31776 = w31784 & w31817;
	assign w31733 = w31776 ^ w31777;
	assign w31761 = w31776 ^ w44702;
	assign w31727 = w31772 ^ w31761;
	assign w31724 = ~w31727;
	assign w31721 = w31777 ^ w31761;
	assign w31737 = w31776 ^ w31779;
	assign w31734 = ~w31737;
	assign w31835 = w31734 ^ w31735;
	assign w31785 = w44704 ^ w31763;
	assign w31783 = w31785 & w31822;
	assign w31774 = w31785 & w31826;
	assign w31750 = w31774 ^ w31749;
	assign w31754 = w31782 ^ w31750;
	assign w31759 = w31783 ^ w31754;
	assign w48893 = w44702 ^ w31759;
	assign w31834 = w31759 ^ w31733;
	assign w31723 = w31781 ^ w31754;
	assign w48892 = w31722 ^ w31723;
	assign w48894 = w31750 ^ w31721;
	assign w7146 = w48890 ^ w48894;
	assign w7177 = w48889 ^ w48893;
	assign w7186 = w48888 ^ w48892;
	assign w44703 = w31781 ^ w31783;
	assign w31739 = w44703 ^ w31736;
	assign w31836 = w31738 ^ w31739;
	assign w31726 = w31730 ^ w44703;
	assign w31729 = w31768 ^ w31726;
	assign w31833 = w31728 ^ w31729;
	assign w31725 = w31749 ^ w31726;
	assign w48891 = w31724 ^ w31725;
	assign w7196 = w48887 ^ w48891;
	assign w7009 = ~w7196;
	assign w45734 = ~w31833;
	assign w7171 = w45561 ^ w45734;
	assign w7006 = w7171 ^ w48893;
	assign w7004 = ~w7006;
	assign w45735 = ~w31834;
	assign w6996 = w7146 ^ w45735;
	assign w7160 = w45554 ^ w45735;
	assign w6999 = w7160 ^ w45734;
	assign w45736 = ~w31835;
	assign w7007 = w7009 ^ w45736;
	assign w7200 = w45555 ^ w45736;
	assign w45737 = ~w31836;
	assign w7208 = w45556 ^ w45737;
	assign w45906 = ~w6665;
	assign w6656 = w45906 ^ w45743;
	assign w6628 = w45906 ^ w45564;
	assign w48613 = w6656 ^ w6657;
	assign w47533 = w48613 ^ w1890;
	assign w48631 = w6627 ^ w6628;
	assign w6625 = w45906 ^ w48695;
	assign w6623 = w6624 ^ w6625;
	assign w48633 = ~w6623;
	assign w47513 = w48633 ^ w1909;
	assign w28502 = w47513 ^ w47514;
	assign w6801 = w47535 ^ w47533;
	assign w6889 = w47536 ^ w47533;
	assign w6884 = w6801 ^ w6807;
	assign w6876 = w6801 ^ w6891;
	assign w6885 = w6889 ^ w6817;
	assign w6882 = w6817 ^ w6884;
	assign w6881 = w6800 ^ w6889;
	assign w6880 = w47540 ^ w6881;
	assign w6763 = w6803 ^ w6801;
	assign w6879 = w6800 ^ w6763;
	assign w6874 = w6881 & w6885;
	assign w6806 = w6874 ^ w6803;
	assign w6873 = w6882 & w6880;
	assign w6869 = w6884 & w6877;
	assign w6890 = w47533 ^ w47539;
	assign w6888 = w47533 ^ w47538;
	assign w6871 = w6890 & w6875;
	assign w6805 = w6871 ^ w6801;
	assign w6868 = w6889 & w6878;
	assign w6804 = w6868 ^ w6802;
	assign w6810 = w6806 ^ w6804;
	assign w6815 = w47533 ^ w6810;
	assign w6867 = w6891 & w6876;
	assign w6776 = w6867 ^ w6868;
	assign w6823 = w6776 ^ w6777;
	assign w6822 = w6823 ^ w6805;
	assign w6864 = w6870 ^ w6822;
	assign w47515 = w48631 ^ w1907;
	assign w28525 = w47515 ^ w47513;
	assign w28527 = w47514 ^ w28525;
	assign w28603 = w47510 ^ w28527;
	assign w28600 = w47511 ^ w28527;
	assign w28602 = w28532 ^ w28527;
	assign w28608 = w47515 ^ w28612;
	assign w28606 = w28525 ^ w28614;
	assign w28605 = w47516 ^ w28606;
	assign w28542 = w47515 ^ w47514;
	assign w28607 = w28542 ^ w28609;
	assign w28610 = w28614 ^ w28542;
	assign w28604 = w28525 ^ w28488;
	assign w28615 = w47509 ^ w47515;
	assign w28599 = w28606 & w28610;
	assign w28531 = w28599 ^ w28528;
	assign w28598 = w28607 & w28605;
	assign w28549 = w28592 ^ w28598;
	assign w28596 = w28615 & w28600;
	assign w28530 = w28596 ^ w28526;
	assign w28595 = w28612 & w28608;
	assign w28594 = w28609 & w28602;
	assign w28593 = w28614 & w28603;
	assign w28529 = w28593 ^ w28527;
	assign w28535 = w28531 ^ w28529;
	assign w28540 = w47509 ^ w28535;
	assign w28590 = w28549 ^ w28540;
	assign w28501 = w28592 ^ w28593;
	assign w28548 = w28501 ^ w28502;
	assign w28547 = w28548 ^ w28530;
	assign w28589 = w28595 ^ w28547;
	assign w28591 = w28613 & w28604;
	assign w28586 = w28590 & w28589;
	assign w6824 = w6867 ^ w6873;
	assign w6865 = w6824 ^ w6815;
	assign w6861 = w6865 & w6864;
	assign w44563 = w28591 ^ w28594;
	assign w28504 = w28530 ^ w44563;
	assign w28588 = w28504 ^ w28529;
	assign w28585 = w28586 ^ w28588;
	assign w28544 = w28592 ^ w44563;
	assign w28500 = w28595 ^ w28544;
	assign w28582 = w47515 ^ w28500;
	assign w44566 = w28591 ^ w28597;
	assign w28503 = w28535 ^ w44566;
	assign w28546 = w47511 ^ w28503;
	assign w28581 = w28586 ^ w28546;
	assign w28580 = w28581 & w28582;
	assign w28578 = w28586 ^ w28580;
	assign w28499 = w28580 ^ w28544;
	assign w28498 = w28580 ^ w28597;
	assign w28493 = w28498 ^ w28594;
	assign w28577 = w28588 & w28578;
	assign w28575 = w28577 ^ w28585;
	assign w44565 = w28577 ^ w28595;
	assign w28569 = w44565 ^ w28547;
	assign w28558 = w28569 & w28610;
	assign w28567 = w28569 & w28606;
	assign w28536 = w47515 ^ w44565;
	assign w28576 = w28536 ^ w28499;
	assign w28566 = w28576 & w28605;
	assign w28557 = w28576 & w28607;
	assign w28579 = w28580 ^ w28588;
	assign w28565 = w28579 & w47516;
	assign w28556 = w28579 & w28611;
	assign w28541 = w44566 ^ w28526;
	assign w28587 = w28549 ^ w28541;
	assign w28584 = w28587 & w28585;
	assign w28583 = w28584 ^ w28546;
	assign w28495 = w28584 ^ w28596;
	assign w28491 = w28495 ^ w28531;
	assign w28494 = w47509 ^ w28491;
	assign w28571 = w28493 ^ w28494;
	assign w28492 = w28584 ^ w28540;
	assign w28490 = w47511 ^ w28491;
	assign w28574 = w28583 & w28575;
	assign w28539 = w28574 ^ w28549;
	assign w28573 = w28539 ^ w28541;
	assign w28497 = w28574 ^ w28598;
	assign w28489 = w28536 ^ w28497;
	assign w28496 = w28526 ^ w28489;
	assign w28572 = w28493 ^ w28496;
	assign w28570 = w28539 ^ w28492;
	assign w28568 = w28489 ^ w28490;
	assign w28564 = w28570 & w28600;
	assign w28563 = w28573 & w28612;
	assign w28562 = w28583 & w28602;
	assign w28506 = w28562 ^ w28563;
	assign w28561 = w28571 & w28603;
	assign w28560 = w28568 & w28601;
	assign w28521 = w28560 ^ w28563;
	assign w28518 = ~w28521;
	assign w28517 = w28560 ^ w28561;
	assign w28559 = w28572 & w28604;
	assign w28555 = w28570 & w28615;
	assign w28537 = w28555 ^ w28559;
	assign w28522 = w28564 ^ w28555;
	assign w28515 = ~w28537;
	assign w28554 = w28573 & w28608;
	assign w28524 = w28562 ^ w28554;
	assign w28553 = w28583 & w28609;
	assign w28514 = w28515 ^ w28553;
	assign w28552 = w28571 & w28614;
	assign w28551 = w28568 & w28616;
	assign w28550 = w28572 & w28613;
	assign w28516 = w28561 ^ w28550;
	assign w28512 = ~w28516;
	assign w44564 = w28551 ^ w28552;
	assign w28533 = w28557 ^ w44564;
	assign w28534 = w28558 ^ w28533;
	assign w28538 = w28566 ^ w28534;
	assign w28507 = w28565 ^ w28538;
	assign w48909 = w28506 ^ w28507;
	assign w28543 = w28567 ^ w28538;
	assign w28618 = w28543 ^ w28517;
	assign w28520 = w28524 ^ w44564;
	assign w28519 = w28515 ^ w28520;
	assign w28619 = w28518 ^ w28519;
	assign w44567 = w28563 ^ w28564;
	assign w48910 = w44567 ^ w28543;
	assign w7161 = w48906 ^ w48910;
	assign w28545 = w28560 ^ w44567;
	assign w28511 = w28556 ^ w28545;
	assign w28508 = ~w28511;
	assign w28505 = w28561 ^ w28545;
	assign w48911 = w28534 ^ w28505;
	assign w7144 = w48907 ^ w48911;
	assign w6951 = w7144 ^ w48909;
	assign w7216 = w6951 ^ w6952;
	assign w44568 = w28565 ^ w28567;
	assign w28523 = w44568 ^ w28520;
	assign w28620 = w28522 ^ w28523;
	assign w28510 = w28514 ^ w44568;
	assign w28513 = w28552 ^ w28510;
	assign w28617 = w28512 ^ w28513;
	assign w28509 = w28533 ^ w28510;
	assign w48908 = w28508 ^ w28509;
	assign w6913 = w48909 ^ w48908;
	assign w7162 = w48904 ^ w48908;
	assign w6866 = w6888 & w6879;
	assign w43786 = w6866 ^ w6872;
	assign w6778 = w6810 ^ w43786;
	assign w6821 = w47535 ^ w6778;
	assign w6856 = w6861 ^ w6821;
	assign w6816 = w43786 ^ w6801;
	assign w6862 = w6824 ^ w6816;
	assign w43787 = w6866 ^ w6869;
	assign w6819 = w6867 ^ w43787;
	assign w6775 = w6870 ^ w6819;
	assign w6857 = w47539 ^ w6775;
	assign w6855 = w6856 & w6857;
	assign w6774 = w6855 ^ w6819;
	assign w6853 = w6861 ^ w6855;
	assign w6773 = w6855 ^ w6872;
	assign w6768 = w6773 ^ w6869;
	assign w6779 = w6805 ^ w43787;
	assign w6863 = w6779 ^ w6804;
	assign w6860 = w6861 ^ w6863;
	assign w6854 = w6855 ^ w6863;
	assign w6831 = w6854 & w6886;
	assign w6859 = w6862 & w6860;
	assign w6770 = w6859 ^ w6871;
	assign w6766 = w6770 ^ w6806;
	assign w6769 = w47533 ^ w6766;
	assign w6767 = w6859 ^ w6815;
	assign w6765 = w47535 ^ w6766;
	assign w6840 = w6854 & w47540;
	assign w6852 = w6863 & w6853;
	assign w6850 = w6852 ^ w6860;
	assign w43791 = w6852 ^ w6870;
	assign w6844 = w43791 ^ w6822;
	assign w6833 = w6844 & w6885;
	assign w6842 = w6844 & w6881;
	assign w43790 = w6840 ^ w6842;
	assign w6811 = w47539 ^ w43791;
	assign w6851 = w6811 ^ w6774;
	assign w6841 = w6851 & w6880;
	assign w6832 = w6851 & w6882;
	assign w6858 = w6859 ^ w6821;
	assign w6828 = w6858 & w6884;
	assign w6837 = w6858 & w6877;
	assign w6846 = w6768 ^ w6769;
	assign w6827 = w6846 & w6889;
	assign w6836 = w6846 & w6878;
	assign w6849 = w6858 & w6850;
	assign w6814 = w6849 ^ w6824;
	assign w6848 = w6814 ^ w6816;
	assign w6845 = w6814 ^ w6767;
	assign w6839 = w6845 & w6875;
	assign w6830 = w6845 & w6890;
	assign w6797 = w6839 ^ w6830;
	assign w6829 = w6848 & w6883;
	assign w6799 = w6837 ^ w6829;
	assign w6838 = w6848 & w6887;
	assign w6781 = w6837 ^ w6838;
	assign w43789 = w6838 ^ w6839;
	assign w6772 = w6849 ^ w6873;
	assign w6764 = w6811 ^ w6772;
	assign w6771 = w6801 ^ w6764;
	assign w6847 = w6768 ^ w6771;
	assign w6834 = w6847 & w6879;
	assign w6812 = w6830 ^ w6834;
	assign w6790 = ~w6812;
	assign w6789 = w6790 ^ w6828;
	assign w6785 = w6789 ^ w43790;
	assign w6825 = w6847 & w6888;
	assign w6791 = w6836 ^ w6825;
	assign w6787 = ~w6791;
	assign w6843 = w6764 ^ w6765;
	assign w6826 = w6843 & w6891;
	assign w6835 = w6843 & w6876;
	assign w6792 = w6835 ^ w6836;
	assign w6796 = w6835 ^ w6838;
	assign w6820 = w6835 ^ w43789;
	assign w6780 = w6836 ^ w6820;
	assign w6793 = ~w6796;
	assign w6788 = w6827 ^ w6785;
	assign w6892 = w6787 ^ w6788;
	assign w43788 = w6826 ^ w6827;
	assign w6808 = w6832 ^ w43788;
	assign w6809 = w6833 ^ w6808;
	assign w48879 = w6809 ^ w6780;
	assign w7154 = w48879 ^ w48894;
	assign w6927 = w7154 ^ w48892;
	assign w6923 = ~w7154;
	assign w6921 = w6923 ^ w45737;
	assign w6924 = w6923 ^ w48891;
	assign w7010 = w7208 ^ w7154;
	assign w6813 = w6841 ^ w6809;
	assign w6818 = w6842 ^ w6813;
	assign w48878 = w43789 ^ w6818;
	assign w6784 = w6808 ^ w6785;
	assign w6893 = w6818 ^ w6792;
	assign w6795 = w6799 ^ w43788;
	assign w6794 = w6790 ^ w6795;
	assign w6798 = w43790 ^ w6795;
	assign w6894 = w6793 ^ w6794;
	assign w6895 = w6797 ^ w6798;
	assign w6786 = w6831 ^ w6820;
	assign w6783 = ~w6786;
	assign w48876 = w6783 ^ w6784;
	assign w6782 = w6840 ^ w6813;
	assign w48877 = w6781 ^ w6782;
	assign w45193 = ~w6893;
	assign w45194 = ~w6894;
	assign w45195 = ~w6895;
	assign w45196 = ~w6892;
	assign w45646 = ~w28617;
	assign w45647 = ~w28618;
	assign w7167 = w45451 ^ w45647;
	assign w45648 = ~w28619;
	assign w7174 = w45452 ^ w45648;
	assign w45649 = ~w28620;
	assign w7194 = w45453 ^ w45649;
	assign w45907 = ~w6672;
	assign w6596 = w45907 ^ w48657;
	assign w6617 = w45907 ^ w48640;
	assign w48522 = w6616 ^ w6617;
	assign w47624 = w48522 ^ w1990;
	assign w14008 = w47624 ^ w47621;
	assign w14010 = w47626 ^ w47624;
	assign w13995 = w13920 ^ w14010;
	assign w13986 = w14010 & w13995;
	assign w13922 = w47624 ^ w47622;
	assign w13882 = w13922 ^ w13920;
	assign w13881 = w13922 ^ w47623;
	assign w14005 = w47628 ^ w13881;
	assign w13991 = w47628 & w14005;
	assign w48533 = w6596 ^ w6597;
	assign w47613 = w48533 ^ w2001;
	assign w20620 = w47615 ^ w47613;
	assign w20695 = w20620 ^ w20710;
	assign w20708 = w47616 ^ w47613;
	assign w20704 = w20708 ^ w20636;
	assign w20703 = w20620 ^ w20626;
	assign w20701 = w20636 ^ w20703;
	assign w20700 = w20619 ^ w20708;
	assign w20699 = w47620 ^ w20700;
	assign w20582 = w20622 ^ w20620;
	assign w20698 = w20619 ^ w20582;
	assign w20709 = w47613 ^ w47619;
	assign w20707 = w47613 ^ w47618;
	assign w20693 = w20700 & w20704;
	assign w20625 = w20693 ^ w20622;
	assign w20692 = w20701 & w20699;
	assign w20690 = w20709 & w20694;
	assign w20624 = w20690 ^ w20620;
	assign w20688 = w20703 & w20696;
	assign w20687 = w20708 & w20697;
	assign w20623 = w20687 ^ w20621;
	assign w20629 = w20625 ^ w20623;
	assign w20634 = w47613 ^ w20629;
	assign w20686 = w20710 & w20695;
	assign w20643 = w20686 ^ w20692;
	assign w20684 = w20643 ^ w20634;
	assign w20595 = w20686 ^ w20687;
	assign w20642 = w20595 ^ w20596;
	assign w20641 = w20642 ^ w20624;
	assign w20683 = w20689 ^ w20641;
	assign w20685 = w20707 & w20698;
	assign w20680 = w20684 & w20683;
	assign w6460 = w45907 ^ w45192;
	assign w6742 = w6460 ^ w6461;
	assign w48519 = w6742 ^ w6734;
	assign w47627 = w48519 ^ w1987;
	assign w14002 = w47627 ^ w14006;
	assign w13936 = w47627 ^ w47626;
	assign w14009 = w47621 ^ w47627;
	assign w13919 = w47627 ^ w47625;
	assign w14000 = w13919 ^ w14008;
	assign w13999 = w47628 ^ w14000;
	assign w13998 = w13919 ^ w13882;
	assign w13985 = w14007 & w13998;
	assign w13989 = w14006 & w14002;
	assign w14004 = w14008 ^ w13936;
	assign w13993 = w14000 & w14004;
	assign w13925 = w13993 ^ w13922;
	assign w14001 = w13936 ^ w14003;
	assign w13992 = w14001 & w13999;
	assign w13921 = w47626 ^ w13919;
	assign w13997 = w47622 ^ w13921;
	assign w13994 = w47623 ^ w13921;
	assign w13990 = w14009 & w13994;
	assign w13924 = w13990 ^ w13920;
	assign w13996 = w13926 ^ w13921;
	assign w13943 = w13986 ^ w13992;
	assign w13988 = w14003 & w13996;
	assign w43953 = w13985 ^ w13991;
	assign w13935 = w43953 ^ w13920;
	assign w13981 = w13943 ^ w13935;
	assign w43954 = w13985 ^ w13988;
	assign w13938 = w13986 ^ w43954;
	assign w13894 = w13989 ^ w13938;
	assign w13976 = w47627 ^ w13894;
	assign w13898 = w13924 ^ w43954;
	assign w44233 = w20685 ^ w20691;
	assign w20635 = w44233 ^ w20620;
	assign w20681 = w20643 ^ w20635;
	assign w20597 = w20629 ^ w44233;
	assign w20640 = w47615 ^ w20597;
	assign w20675 = w20680 ^ w20640;
	assign w44234 = w20685 ^ w20688;
	assign w20638 = w20686 ^ w44234;
	assign w20594 = w20689 ^ w20638;
	assign w20676 = w47619 ^ w20594;
	assign w20674 = w20675 & w20676;
	assign w20593 = w20674 ^ w20638;
	assign w20592 = w20674 ^ w20691;
	assign w20587 = w20592 ^ w20688;
	assign w20672 = w20680 ^ w20674;
	assign w20598 = w20624 ^ w44234;
	assign w20682 = w20598 ^ w20623;
	assign w20673 = w20674 ^ w20682;
	assign w20679 = w20680 ^ w20682;
	assign w20678 = w20681 & w20679;
	assign w20677 = w20678 ^ w20640;
	assign w20589 = w20678 ^ w20690;
	assign w20585 = w20589 ^ w20625;
	assign w20588 = w47613 ^ w20585;
	assign w20665 = w20587 ^ w20588;
	assign w20586 = w20678 ^ w20634;
	assign w20584 = w47615 ^ w20585;
	assign w20671 = w20682 & w20672;
	assign w20669 = w20671 ^ w20679;
	assign w20668 = w20677 & w20669;
	assign w20633 = w20668 ^ w20643;
	assign w20667 = w20633 ^ w20635;
	assign w20591 = w20668 ^ w20692;
	assign w20664 = w20633 ^ w20586;
	assign w20659 = w20673 & w47620;
	assign w20658 = w20664 & w20694;
	assign w20657 = w20667 & w20706;
	assign w20656 = w20677 & w20696;
	assign w20600 = w20656 ^ w20657;
	assign w20655 = w20665 & w20697;
	assign w20650 = w20673 & w20705;
	assign w20649 = w20664 & w20709;
	assign w20616 = w20658 ^ w20649;
	assign w20648 = w20667 & w20702;
	assign w20618 = w20656 ^ w20648;
	assign w20647 = w20677 & w20703;
	assign w20646 = w20665 & w20708;
	assign w44235 = w20657 ^ w20658;
	assign w44237 = w20671 ^ w20689;
	assign w20630 = w47619 ^ w44237;
	assign w20670 = w20630 ^ w20593;
	assign w20651 = w20670 & w20701;
	assign w20660 = w20670 & w20699;
	assign w20583 = w20630 ^ w20591;
	assign w20590 = w20620 ^ w20583;
	assign w20666 = w20587 ^ w20590;
	assign w20653 = w20666 & w20698;
	assign w20631 = w20649 ^ w20653;
	assign w20609 = ~w20631;
	assign w20608 = w20609 ^ w20647;
	assign w20662 = w20583 ^ w20584;
	assign w20645 = w20662 & w20710;
	assign w20644 = w20666 & w20707;
	assign w20610 = w20655 ^ w20644;
	assign w20606 = ~w20610;
	assign w43556 = w20645 ^ w20646;
	assign w20627 = w20651 ^ w43556;
	assign w20614 = w20618 ^ w43556;
	assign w20613 = w20609 ^ w20614;
	assign w20654 = w20662 & w20695;
	assign w20611 = w20654 ^ w20655;
	assign w20639 = w20654 ^ w44235;
	assign w20605 = w20650 ^ w20639;
	assign w20602 = ~w20605;
	assign w20599 = w20655 ^ w20639;
	assign w20615 = w20654 ^ w20657;
	assign w20612 = ~w20615;
	assign w20713 = w20612 ^ w20613;
	assign w20663 = w44237 ^ w20641;
	assign w20661 = w20663 & w20700;
	assign w20652 = w20663 & w20704;
	assign w20628 = w20652 ^ w20627;
	assign w20632 = w20660 ^ w20628;
	assign w20637 = w20661 ^ w20632;
	assign w48870 = w44235 ^ w20637;
	assign w20712 = w20637 ^ w20611;
	assign w20601 = w20659 ^ w20632;
	assign w48869 = w20600 ^ w20601;
	assign w48871 = w20628 ^ w20599;
	assign w7017 = ~w48870;
	assign w7032 = w7017 ^ w48866;
	assign w48764 = w7031 ^ w7032;
	assign w6919 = w48869 ^ w6907;
	assign w47455 = w48764 ^ w1426;
	assign w7155 = w48867 ^ w48871;
	assign w6916 = w7155 ^ w48873;
	assign w6920 = ~w7155;
	assign w6918 = w6920 ^ w48874;
	assign w6914 = w7155 ^ w45740;
	assign w7173 = w48869 ^ w48873;
	assign w7015 = w7018 ^ w7173;
	assign w48746 = w7235 ^ w7173;
	assign w47473 = w48746 ^ w1408;
	assign w7147 = w48871 ^ w48875;
	assign w7056 = w7166 ^ w7147;
	assign w48750 = w48867 ^ w7056;
	assign w7027 = w7188 ^ w7147;
	assign w7023 = w7147 ^ w48869;
	assign w7038 = w7147 ^ w45272;
	assign w7016 = w7147 ^ w7017;
	assign w48771 = w7015 ^ w7016;
	assign w47448 = w48771 ^ w1433;
	assign w7168 = w48870 ^ w48874;
	assign w7042 = w7044 ^ w7168;
	assign w7014 = w7172 ^ w7168;
	assign w48747 = w7234 ^ w7168;
	assign w47472 = w48747 ^ w1409;
	assign w48758 = w7038 ^ w7039;
	assign w47461 = w48758 ^ w1420;
	assign w7045 = w7036 ^ w7173;
	assign w7037 = w7188 ^ w7155;
	assign w48759 = w45741 ^ w7037;
	assign w47460 = w48759 ^ w1421;
	assign w47469 = w48750 ^ w1412;
	assign w19904 = w47472 ^ w47469;
	assign w44236 = w20659 ^ w20661;
	assign w20617 = w44236 ^ w20614;
	assign w20714 = w20616 ^ w20617;
	assign w20604 = w20608 ^ w44236;
	assign w20607 = w20646 ^ w20604;
	assign w20711 = w20606 ^ w20607;
	assign w20603 = w20627 ^ w20604;
	assign w48868 = w20602 ^ w20603;
	assign w6917 = w48868 ^ w48864;
	assign w7230 = w6916 ^ w6917;
	assign w48762 = w7230 ^ w7180;
	assign w47457 = w48762 ^ w1424;
	assign w7178 = w48868 ^ w48872;
	assign w7061 = w7178 ^ w45740;
	assign w7022 = w7180 ^ w7178;
	assign w48770 = w7022 ^ w7023;
	assign w47449 = w48770 ^ w1432;
	assign w7047 = w7187 ^ w7178;
	assign w48753 = w48859 ^ w7047;
	assign w47466 = w48753 ^ w1415;
	assign w34241 = w47461 ^ w47466;
	assign w48745 = w7061 ^ w7062;
	assign w47474 = w48745 ^ w1407;
	assign w19906 = w47474 ^ w47472;
	assign w19792 = w47473 ^ w47474;
	assign w19903 = w47469 ^ w47474;
	assign w13987 = w14008 & w13997;
	assign w13923 = w13987 ^ w13921;
	assign w13929 = w13925 ^ w13923;
	assign w13934 = w47621 ^ w13929;
	assign w13982 = w13898 ^ w13923;
	assign w13897 = w13929 ^ w43953;
	assign w13984 = w13943 ^ w13934;
	assign w13940 = w47623 ^ w13897;
	assign w13895 = w13986 ^ w13987;
	assign w13942 = w13895 ^ w13896;
	assign w13941 = w13942 ^ w13924;
	assign w13983 = w13989 ^ w13941;
	assign w13980 = w13984 & w13983;
	assign w13975 = w13980 ^ w13940;
	assign w13974 = w13975 & w13976;
	assign w13973 = w13974 ^ w13982;
	assign w13892 = w13974 ^ w13991;
	assign w13887 = w13892 ^ w13988;
	assign w13950 = w13973 & w14005;
	assign w13959 = w13973 & w47628;
	assign w13979 = w13980 ^ w13982;
	assign w13978 = w13981 & w13979;
	assign w13977 = w13978 ^ w13940;
	assign w13889 = w13978 ^ w13990;
	assign w13886 = w13978 ^ w13934;
	assign w13972 = w13980 ^ w13974;
	assign w13893 = w13974 ^ w13938;
	assign w13885 = w13889 ^ w13925;
	assign w13888 = w47621 ^ w13885;
	assign w13965 = w13887 ^ w13888;
	assign w13884 = w47623 ^ w13885;
	assign w13955 = w13965 & w13997;
	assign w13947 = w13977 & w14003;
	assign w13956 = w13977 & w13996;
	assign w13971 = w13982 & w13972;
	assign w13969 = w13971 ^ w13979;
	assign w13968 = w13977 & w13969;
	assign w13933 = w13968 ^ w13943;
	assign w13967 = w13933 ^ w13935;
	assign w13891 = w13968 ^ w13992;
	assign w13964 = w13933 ^ w13886;
	assign w13949 = w13964 & w14009;
	assign w13958 = w13964 & w13994;
	assign w13916 = w13958 ^ w13949;
	assign w13948 = w13967 & w14002;
	assign w13918 = w13956 ^ w13948;
	assign w13957 = w13967 & w14006;
	assign w13900 = w13956 ^ w13957;
	assign w43955 = w13957 ^ w13958;
	assign w43957 = w13971 ^ w13989;
	assign w13930 = w47627 ^ w43957;
	assign w13883 = w13930 ^ w13891;
	assign w13962 = w13883 ^ w13884;
	assign w13945 = w13962 & w14010;
	assign w13890 = w13920 ^ w13883;
	assign w13966 = w13887 ^ w13890;
	assign w13944 = w13966 & w14007;
	assign w13910 = w13955 ^ w13944;
	assign w13906 = ~w13910;
	assign w13953 = w13966 & w13998;
	assign w13931 = w13949 ^ w13953;
	assign w13909 = ~w13931;
	assign w13908 = w13909 ^ w13947;
	assign w13970 = w13930 ^ w13893;
	assign w13951 = w13970 & w14001;
	assign w13960 = w13970 & w13999;
	assign w13963 = w43957 ^ w13941;
	assign w13952 = w13963 & w14004;
	assign w13961 = w13963 & w14000;
	assign w43956 = w13959 ^ w13961;
	assign w13904 = w13908 ^ w43956;
	assign w13954 = w13962 & w13995;
	assign w13939 = w13954 ^ w43955;
	assign w13899 = w13955 ^ w13939;
	assign w13905 = w13950 ^ w13939;
	assign w13902 = ~w13905;
	assign w13915 = w13954 ^ w13957;
	assign w13912 = ~w13915;
	assign w13911 = w13954 ^ w13955;
	assign w7229 = w6918 ^ w6919;
	assign w48763 = w7229 ^ w7176;
	assign w47456 = w48763 ^ w1425;
	assign w13946 = w13965 & w14008;
	assign w13907 = w13946 ^ w13904;
	assign w14011 = w13906 ^ w13907;
	assign w6974 = w45561 ^ w14011;
	assign w7005 = w14011 ^ w48878;
	assign w48780 = w7004 ^ w7005;
	assign w47439 = w48780 ^ w1378;
	assign w48884 = ~w14011;
	assign w7182 = w45196 ^ w48884;
	assign w6985 = w7182 ^ w7160;
	assign w6976 = w7182 ^ w45734;
	assign w48789 = w45193 ^ w6985;
	assign w6958 = w7182 ^ w7177;
	assign w48804 = w45561 ^ w6958;
	assign w47430 = w48789 ^ w1387;
	assign w47415 = w48804 ^ w1402;
	assign w43536 = w13945 ^ w13946;
	assign w13914 = w13918 ^ w43536;
	assign w13913 = w13909 ^ w13914;
	assign w13917 = w43956 ^ w13914;
	assign w14013 = w13912 ^ w13913;
	assign w6922 = w14013 ^ w45195;
	assign w7228 = w6921 ^ w6922;
	assign w48776 = w7228 ^ w7200;
	assign w47443 = w48776 ^ w1374;
	assign w6979 = w45555 ^ w14013;
	assign w14014 = w13916 ^ w13917;
	assign w48880 = ~w14013;
	assign w7211 = w45194 ^ w48880;
	assign w6991 = w7211 ^ w7196;
	assign w48785 = w48876 ^ w6991;
	assign w47434 = w48785 ^ w1383;
	assign w6969 = w7211 ^ w7208;
	assign w6967 = ~w6969;
	assign w13927 = w13951 ^ w43536;
	assign w13928 = w13952 ^ w13927;
	assign w48886 = w13928 ^ w13899;
	assign w13903 = w13927 ^ w13904;
	assign w48881 = w13902 ^ w13903;
	assign w6997 = w48886 ^ w45193;
	assign w48782 = w6996 ^ w6997;
	assign w6933 = ~w48881;
	assign w7008 = w6933 ^ w45194;
	assign w48777 = w7007 ^ w7008;
	assign w47437 = w48782 ^ w1380;
	assign w25042 = w47439 ^ w47437;
	assign w25131 = w47437 ^ w47443;
	assign w47442 = w48777 ^ w1375;
	assign w25058 = w47443 ^ w47442;
	assign w25129 = w47437 ^ w47442;
	assign w7149 = w48879 ^ w48886;
	assign w6995 = w7208 ^ w7149;
	assign w48783 = w45195 ^ w6995;
	assign w6956 = w7160 ^ w7149;
	assign w48806 = w48890 ^ w6956;
	assign w47436 = w48783 ^ w1381;
	assign w13390 = w47436 ^ w47430;
	assign w47413 = w48806 ^ w1404;
	assign w28392 = w47415 ^ w47413;
	assign w7153 = w48886 ^ w48890;
	assign w6934 = ~w7153;
	assign w6931 = w6934 ^ w48892;
	assign w6935 = w6934 ^ w48893;
	assign w6929 = w7153 ^ w45736;
	assign w7204 = w48876 ^ w48881;
	assign w6965 = w7204 ^ w7200;
	assign w6980 = ~w7204;
	assign w6978 = w6980 ^ w48891;
	assign w48793 = w6978 ^ w6979;
	assign w48801 = w48887 ^ w6965;
	assign w6989 = w6980 ^ w7186;
	assign w47418 = w48801 ^ w1399;
	assign w28479 = w47413 ^ w47418;
	assign w47426 = w48793 ^ w1391;
	assign w13932 = w13960 ^ w13928;
	assign w13901 = w13959 ^ w13932;
	assign w13937 = w13961 ^ w13932;
	assign w48883 = w43955 ^ w13937;
	assign w14012 = w13937 ^ w13911;
	assign w48882 = w13900 ^ w13901;
	assign w6928 = w48883 ^ w48877;
	assign w6977 = w48889 ^ w48883;
	assign w6926 = ~w48882;
	assign w48796 = w6976 ^ w6977;
	assign w7226 = w6927 ^ w6928;
	assign w6936 = w48888 ^ w6926;
	assign w7223 = w6935 ^ w6936;
	assign w6925 = w6926 ^ w48876;
	assign w7227 = w6924 ^ w6925;
	assign w7000 = w14012 ^ w45196;
	assign w6998 = w6999 ^ w7000;
	assign w48781 = ~w6998;
	assign w6972 = w45554 ^ w14012;
	assign w47438 = w48781 ^ w1379;
	assign w47423 = w48796 ^ w1394;
	assign w48885 = ~w14012;
	assign w48778 = w7227 ^ w7186;
	assign w47441 = w48778 ^ w1376;
	assign w25041 = w47443 ^ w47441;
	assign w25043 = w47442 ^ w25041;
	assign w25119 = w47438 ^ w25043;
	assign w25116 = w47439 ^ w25043;
	assign w25018 = w47441 ^ w47442;
	assign w25112 = w25131 & w25116;
	assign w25046 = w25112 ^ w25042;
	assign w48779 = w7226 ^ w7177;
	assign w47440 = w48779 ^ w1377;
	assign w25044 = w47440 ^ w47438;
	assign w25130 = w47440 ^ w47437;
	assign w25126 = w25130 ^ w25058;
	assign w25122 = w25041 ^ w25130;
	assign w25132 = w47442 ^ w47440;
	assign w25117 = w25042 ^ w25132;
	assign w25004 = w25044 ^ w25042;
	assign w25120 = w25041 ^ w25004;
	assign w25003 = w25044 ^ w47439;
	assign w25115 = w25122 & w25126;
	assign w25047 = w25115 ^ w25044;
	assign w25109 = w25130 & w25119;
	assign w25045 = w25109 ^ w25043;
	assign w25051 = w25047 ^ w25045;
	assign w25056 = w47437 ^ w25051;
	assign w25108 = w25132 & w25117;
	assign w25017 = w25108 ^ w25109;
	assign w25064 = w25017 ^ w25018;
	assign w25063 = w25064 ^ w25046;
	assign w25107 = w25129 & w25120;
	assign w7175 = w45193 ^ w48885;
	assign w6984 = w7175 ^ w7146;
	assign w48790 = w48879 ^ w6984;
	assign w6975 = w7175 ^ w45735;
	assign w6973 = ~w6975;
	assign w6957 = w7175 ^ w7171;
	assign w48805 = w45554 ^ w6957;
	assign w47429 = w48790 ^ w1388;
	assign w13471 = w47429 ^ w47434;
	assign w47414 = w48805 ^ w1403;
	assign w7197 = w48877 ^ w48882;
	assign w6964 = ~w7197;
	assign w6962 = w6964 ^ w7196;
	assign w6987 = w6964 ^ w7177;
	assign w7189 = w48878 ^ w48883;
	assign w6986 = w7189 ^ w7171;
	assign w48788 = w45196 ^ w6986;
	assign w6961 = ~w7189;
	assign w6959 = w6961 ^ w7186;
	assign w47431 = w48788 ^ w1386;
	assign w13470 = w47431 ^ w13390;
	assign w13384 = w47431 ^ w47429;
	assign w13467 = w13384 ^ w13390;
	assign w48795 = w7223 ^ w7189;
	assign w47424 = w48795 ^ w1393;
	assign w19638 = w47426 ^ w47424;
	assign w48797 = w6973 ^ w6974;
	assign w47422 = w48797 ^ w1395;
	assign w19550 = w47424 ^ w47422;
	assign w19509 = w19550 ^ w47423;
	assign w6932 = w48887 ^ w6933;
	assign w7224 = w6931 ^ w6932;
	assign w48794 = w7224 ^ w7197;
	assign w47425 = w48794 ^ w1392;
	assign w19524 = w47425 ^ w47426;
	assign w45274 = ~w14014;
	assign w6930 = w45556 ^ w45274;
	assign w7225 = w6929 ^ w6930;
	assign w48775 = w45274 ^ w7010;
	assign w47444 = w48775 ^ w1373;
	assign w25121 = w47444 ^ w25122;
	assign w25048 = w47444 ^ w47438;
	assign w25118 = w25048 ^ w25043;
	assign w25125 = w25042 ^ w25048;
	assign w25123 = w25058 ^ w25125;
	assign w25128 = w47439 ^ w25048;
	assign w25124 = w47443 ^ w25128;
	assign w25127 = w47444 ^ w25003;
	assign w25114 = w25123 & w25121;
	assign w25065 = w25108 ^ w25114;
	assign w25106 = w25065 ^ w25056;
	assign w25113 = w47444 & w25127;
	assign w25111 = w25128 & w25124;
	assign w25105 = w25111 ^ w25063;
	assign w25110 = w25125 & w25118;
	assign w25102 = w25106 & w25105;
	assign w48792 = w7225 ^ w7211;
	assign w47427 = w48792 ^ w1390;
	assign w19547 = w47427 ^ w47425;
	assign w19549 = w47426 ^ w19547;
	assign w19625 = w47422 ^ w19549;
	assign w19622 = w47423 ^ w19549;
	assign w19564 = w47427 ^ w47426;
	assign w7212 = w45195 ^ w45274;
	assign w6981 = w7212 ^ w7153;
	assign w48791 = w45737 ^ w6981;
	assign w6970 = w7212 ^ w7146;
	assign w48799 = w45556 ^ w6970;
	assign w6993 = w7212 ^ w7200;
	assign w47428 = w48791 ^ w1389;
	assign w19554 = w47428 ^ w47422;
	assign w19624 = w19554 ^ w19549;
	assign w19634 = w47423 ^ w19554;
	assign w19630 = w47427 ^ w19634;
	assign w19633 = w47428 ^ w19509;
	assign w19619 = w47428 & w19633;
	assign w19617 = w19634 & w19630;
	assign w47420 = w48799 ^ w1397;
	assign w28398 = w47420 ^ w47414;
	assign w28475 = w28392 ^ w28398;
	assign w28478 = w47415 ^ w28398;
	assign w44419 = w25107 ^ w25113;
	assign w25057 = w44419 ^ w25042;
	assign w25103 = w25065 ^ w25057;
	assign w25019 = w25051 ^ w44419;
	assign w25062 = w47439 ^ w25019;
	assign w25097 = w25102 ^ w25062;
	assign w44420 = w25107 ^ w25110;
	assign w25060 = w25108 ^ w44420;
	assign w25016 = w25111 ^ w25060;
	assign w25098 = w47443 ^ w25016;
	assign w25096 = w25097 & w25098;
	assign w25015 = w25096 ^ w25060;
	assign w25014 = w25096 ^ w25113;
	assign w25009 = w25014 ^ w25110;
	assign w25094 = w25102 ^ w25096;
	assign w25020 = w25046 ^ w44420;
	assign w25104 = w25020 ^ w25045;
	assign w25095 = w25096 ^ w25104;
	assign w25101 = w25102 ^ w25104;
	assign w25100 = w25103 & w25101;
	assign w25099 = w25100 ^ w25062;
	assign w25011 = w25100 ^ w25112;
	assign w25007 = w25011 ^ w25047;
	assign w25010 = w47437 ^ w25007;
	assign w25087 = w25009 ^ w25010;
	assign w25008 = w25100 ^ w25056;
	assign w25006 = w47439 ^ w25007;
	assign w25093 = w25104 & w25094;
	assign w25091 = w25093 ^ w25101;
	assign w25090 = w25099 & w25091;
	assign w25055 = w25090 ^ w25065;
	assign w25089 = w25055 ^ w25057;
	assign w25013 = w25090 ^ w25114;
	assign w25086 = w25055 ^ w25008;
	assign w25081 = w25095 & w47444;
	assign w25080 = w25086 & w25116;
	assign w25079 = w25089 & w25128;
	assign w25078 = w25099 & w25118;
	assign w25022 = w25078 ^ w25079;
	assign w25077 = w25087 & w25119;
	assign w25072 = w25095 & w25127;
	assign w25071 = w25086 & w25131;
	assign w25038 = w25080 ^ w25071;
	assign w25070 = w25089 & w25124;
	assign w25040 = w25078 ^ w25070;
	assign w25069 = w25099 & w25125;
	assign w25068 = w25087 & w25130;
	assign w44421 = w25079 ^ w25080;
	assign w44423 = w25093 ^ w25111;
	assign w25052 = w47443 ^ w44423;
	assign w25092 = w25052 ^ w25015;
	assign w25073 = w25092 & w25123;
	assign w25082 = w25092 & w25121;
	assign w25005 = w25052 ^ w25013;
	assign w25012 = w25042 ^ w25005;
	assign w25088 = w25009 ^ w25012;
	assign w25075 = w25088 & w25120;
	assign w25053 = w25071 ^ w25075;
	assign w25031 = ~w25053;
	assign w25030 = w25031 ^ w25069;
	assign w25084 = w25005 ^ w25006;
	assign w25067 = w25084 & w25132;
	assign w25066 = w25088 & w25129;
	assign w25032 = w25077 ^ w25066;
	assign w25028 = ~w25032;
	assign w43568 = w25067 ^ w25068;
	assign w25049 = w25073 ^ w43568;
	assign w25036 = w25040 ^ w43568;
	assign w25035 = w25031 ^ w25036;
	assign w25076 = w25084 & w25117;
	assign w25037 = w25076 ^ w25079;
	assign w25034 = ~w25037;
	assign w25135 = w25034 ^ w25035;
	assign w25033 = w25076 ^ w25077;
	assign w25061 = w25076 ^ w44421;
	assign w25021 = w25077 ^ w25061;
	assign w25027 = w25072 ^ w25061;
	assign w25024 = ~w25027;
	assign w25085 = w44423 ^ w25063;
	assign w25083 = w25085 & w25122;
	assign w25074 = w25085 & w25126;
	assign w25050 = w25074 ^ w25049;
	assign w25054 = w25082 ^ w25050;
	assign w25059 = w25083 ^ w25054;
	assign w49062 = w44421 ^ w25059;
	assign w25134 = w25059 ^ w25033;
	assign w25023 = w25081 ^ w25054;
	assign w49061 = w25022 ^ w25023;
	assign w49063 = w25050 ^ w25021;
	assign w44422 = w25081 ^ w25083;
	assign w25039 = w44422 ^ w25036;
	assign w25136 = w25038 ^ w25039;
	assign w25026 = w25030 ^ w44422;
	assign w25029 = w25068 ^ w25026;
	assign w25133 = w25028 ^ w25029;
	assign w25025 = w25049 ^ w25026;
	assign w49060 = w25024 ^ w25025;
	assign w45462 = ~w20711;
	assign w7029 = w7166 ^ w45462;
	assign w48765 = w7029 ^ w7030;
	assign w48772 = w45462 ^ w7014;
	assign w47447 = w48772 ^ w1434;
	assign w47454 = w48765 ^ w1427;
	assign w19684 = w47456 ^ w47454;
	assign w19688 = w47460 ^ w47454;
	assign w19768 = w47455 ^ w19688;
	assign w19643 = w19684 ^ w47455;
	assign w19767 = w47460 ^ w19643;
	assign w19753 = w47460 & w19767;
	assign w7163 = w45462 ^ w45738;
	assign w7041 = w7176 ^ w7163;
	assign w48756 = w45454 ^ w7041;
	assign w47463 = w48756 ^ w1418;
	assign w34154 = w47463 ^ w47461;
	assign w7059 = w7163 ^ w48874;
	assign w48748 = w7059 ^ w7060;
	assign w47471 = w48748 ^ w1410;
	assign w19816 = w47471 ^ w47469;
	assign w19891 = w19816 ^ w19906;
	assign w19882 = w19906 & w19891;
	assign w45463 = ~w20712;
	assign w7012 = w48871 ^ w45463;
	assign w48774 = w7011 ^ w7012;
	assign w48757 = w45463 ^ w7040;
	assign w47462 = w48757 ^ w1419;
	assign w47445 = w48774 ^ w1436;
	assign w31474 = w47447 ^ w47445;
	assign w31562 = w47448 ^ w47445;
	assign w7165 = w45272 ^ w45463;
	assign w7057 = w7165 ^ w45739;
	assign w48749 = w7057 ^ w7058;
	assign w7028 = w7165 ^ w7148;
	assign w48766 = w48875 ^ w7028;
	assign w7013 = w7165 ^ w7163;
	assign w48773 = w45455 ^ w7013;
	assign w47453 = w48766 ^ w1428;
	assign w19682 = w47455 ^ w47453;
	assign w19770 = w47456 ^ w47453;
	assign w19765 = w19682 ^ w19688;
	assign w19644 = w19684 ^ w19682;
	assign w47470 = w48749 ^ w1411;
	assign w19818 = w47472 ^ w47470;
	assign w19778 = w19818 ^ w19816;
	assign w19777 = w19818 ^ w47471;
	assign w47446 = w48773 ^ w1435;
	assign w31476 = w47448 ^ w47446;
	assign w31436 = w31476 ^ w31474;
	assign w31435 = w31476 ^ w47447;
	assign w45464 = ~w20713;
	assign w7035 = w45464 ^ w13745;
	assign w48761 = w7034 ^ w7035;
	assign w7026 = w7147 ^ w45464;
	assign w47458 = w48761 ^ w1423;
	assign w19772 = w47458 ^ w47456;
	assign w19757 = w19682 ^ w19772;
	assign w19658 = w47457 ^ w47458;
	assign w19769 = w47453 ^ w47458;
	assign w19748 = w19772 & w19757;
	assign w7181 = w45464 ^ w45740;
	assign w7049 = w7188 ^ w7181;
	assign w7024 = w7183 ^ w7181;
	assign w48769 = w48868 ^ w7024;
	assign w47450 = w48769 ^ w1431;
	assign w31564 = w47450 ^ w47448;
	assign w31549 = w31474 ^ w31564;
	assign w31450 = w47449 ^ w47450;
	assign w31561 = w47445 ^ w47450;
	assign w31540 = w31564 & w31549;
	assign w48744 = w7236 ^ w7181;
	assign w47475 = w48744 ^ w1406;
	assign w19815 = w47475 ^ w47473;
	assign w19817 = w47474 ^ w19815;
	assign w19893 = w47470 ^ w19817;
	assign w19890 = w47471 ^ w19817;
	assign w19896 = w19815 ^ w19904;
	assign w19832 = w47475 ^ w47474;
	assign w19900 = w19904 ^ w19832;
	assign w19894 = w19815 ^ w19778;
	assign w19905 = w47469 ^ w47475;
	assign w19889 = w19896 & w19900;
	assign w19821 = w19889 ^ w19818;
	assign w19886 = w19905 & w19890;
	assign w19820 = w19886 ^ w19816;
	assign w19883 = w19904 & w19893;
	assign w19819 = w19883 ^ w19817;
	assign w19825 = w19821 ^ w19819;
	assign w19830 = w47469 ^ w19825;
	assign w19791 = w19882 ^ w19883;
	assign w19838 = w19791 ^ w19792;
	assign w19837 = w19838 ^ w19820;
	assign w19881 = w19903 & w19894;
	assign w45465 = ~w20714;
	assign w48767 = w45465 ^ w7027;
	assign w47452 = w48767 ^ w1429;
	assign w31480 = w47452 ^ w47446;
	assign w31557 = w31474 ^ w31480;
	assign w31560 = w47447 ^ w31480;
	assign w31559 = w47452 ^ w31435;
	assign w31545 = w47452 & w31559;
	assign w7185 = w45465 ^ w45741;
	assign w7025 = w7187 ^ w7185;
	assign w48768 = w7025 ^ w7026;
	assign w47451 = w48768 ^ w1430;
	assign w31473 = w47451 ^ w47449;
	assign w31475 = w47450 ^ w31473;
	assign w31551 = w47446 ^ w31475;
	assign w31548 = w47447 ^ w31475;
	assign w31550 = w31480 ^ w31475;
	assign w31556 = w47451 ^ w31560;
	assign w31554 = w31473 ^ w31562;
	assign w31553 = w47452 ^ w31554;
	assign w31490 = w47451 ^ w47450;
	assign w31555 = w31490 ^ w31557;
	assign w31558 = w31562 ^ w31490;
	assign w31552 = w31473 ^ w31436;
	assign w31563 = w47445 ^ w47451;
	assign w31547 = w31554 & w31558;
	assign w31479 = w31547 ^ w31476;
	assign w31546 = w31555 & w31553;
	assign w31497 = w31540 ^ w31546;
	assign w31544 = w31563 & w31548;
	assign w31478 = w31544 ^ w31474;
	assign w31543 = w31560 & w31556;
	assign w31542 = w31557 & w31550;
	assign w31541 = w31562 & w31551;
	assign w31477 = w31541 ^ w31475;
	assign w31483 = w31479 ^ w31477;
	assign w31488 = w47445 ^ w31483;
	assign w31538 = w31497 ^ w31488;
	assign w31449 = w31540 ^ w31541;
	assign w31496 = w31449 ^ w31450;
	assign w31495 = w31496 ^ w31478;
	assign w31537 = w31543 ^ w31495;
	assign w31539 = w31561 & w31552;
	assign w31534 = w31538 & w31537;
	assign w7063 = w7185 ^ w7157;
	assign w48743 = w45273 ^ w7063;
	assign w7051 = w7185 ^ w7148;
	assign w48751 = w45457 ^ w7051;
	assign w47468 = w48751 ^ w1413;
	assign w34160 = w47468 ^ w47462;
	assign w34237 = w34154 ^ w34160;
	assign w34240 = w47463 ^ w34160;
	assign w47476 = w48743 ^ w1405;
	assign w19895 = w47476 ^ w19896;
	assign w19822 = w47476 ^ w47470;
	assign w19892 = w19822 ^ w19817;
	assign w19899 = w19816 ^ w19822;
	assign w19897 = w19832 ^ w19899;
	assign w19902 = w47471 ^ w19822;
	assign w19898 = w47475 ^ w19902;
	assign w19901 = w47476 ^ w19777;
	assign w19888 = w19897 & w19895;
	assign w19839 = w19882 ^ w19888;
	assign w19880 = w19839 ^ w19830;
	assign w19887 = w47476 & w19901;
	assign w19885 = w19902 & w19898;
	assign w19879 = w19885 ^ w19837;
	assign w19884 = w19899 & w19892;
	assign w19876 = w19880 & w19879;
	assign w44199 = w19881 ^ w19884;
	assign w19794 = w19820 ^ w44199;
	assign w19878 = w19794 ^ w19819;
	assign w19875 = w19876 ^ w19878;
	assign w19834 = w19882 ^ w44199;
	assign w19790 = w19885 ^ w19834;
	assign w19872 = w47475 ^ w19790;
	assign w44202 = w19881 ^ w19887;
	assign w19793 = w19825 ^ w44202;
	assign w19836 = w47471 ^ w19793;
	assign w19871 = w19876 ^ w19836;
	assign w19870 = w19871 & w19872;
	assign w19869 = w19870 ^ w19878;
	assign w19868 = w19876 ^ w19870;
	assign w19789 = w19870 ^ w19834;
	assign w19788 = w19870 ^ w19887;
	assign w19783 = w19788 ^ w19884;
	assign w19867 = w19878 & w19868;
	assign w19865 = w19867 ^ w19875;
	assign w19855 = w19869 & w47476;
	assign w19846 = w19869 & w19901;
	assign w44201 = w19867 ^ w19885;
	assign w19859 = w44201 ^ w19837;
	assign w19857 = w19859 & w19896;
	assign w19848 = w19859 & w19900;
	assign w19826 = w47475 ^ w44201;
	assign w19866 = w19826 ^ w19789;
	assign w19856 = w19866 & w19895;
	assign w19847 = w19866 & w19897;
	assign w19831 = w44202 ^ w19816;
	assign w19877 = w19839 ^ w19831;
	assign w19874 = w19877 & w19875;
	assign w19873 = w19874 ^ w19836;
	assign w19785 = w19874 ^ w19886;
	assign w19781 = w19785 ^ w19821;
	assign w19784 = w47469 ^ w19781;
	assign w19861 = w19783 ^ w19784;
	assign w19782 = w19874 ^ w19830;
	assign w19780 = w47471 ^ w19781;
	assign w19864 = w19873 & w19865;
	assign w19829 = w19864 ^ w19839;
	assign w19863 = w19829 ^ w19831;
	assign w19787 = w19864 ^ w19888;
	assign w19779 = w19826 ^ w19787;
	assign w19786 = w19816 ^ w19779;
	assign w19862 = w19783 ^ w19786;
	assign w19860 = w19829 ^ w19782;
	assign w19858 = w19779 ^ w19780;
	assign w19854 = w19860 & w19890;
	assign w19853 = w19863 & w19902;
	assign w19852 = w19873 & w19892;
	assign w19796 = w19852 ^ w19853;
	assign w19851 = w19861 & w19893;
	assign w19850 = w19858 & w19891;
	assign w19811 = w19850 ^ w19853;
	assign w19808 = ~w19811;
	assign w19807 = w19850 ^ w19851;
	assign w19849 = w19862 & w19894;
	assign w19845 = w19860 & w19905;
	assign w19827 = w19845 ^ w19849;
	assign w19812 = w19854 ^ w19845;
	assign w19805 = ~w19827;
	assign w19844 = w19863 & w19898;
	assign w19814 = w19852 ^ w19844;
	assign w19843 = w19873 & w19899;
	assign w19804 = w19805 ^ w19843;
	assign w19842 = w19861 & w19904;
	assign w19841 = w19858 & w19906;
	assign w19840 = w19862 & w19903;
	assign w19806 = w19851 ^ w19840;
	assign w19802 = ~w19806;
	assign w44200 = w19841 ^ w19842;
	assign w19823 = w19847 ^ w44200;
	assign w19824 = w19848 ^ w19823;
	assign w19828 = w19856 ^ w19824;
	assign w19833 = w19857 ^ w19828;
	assign w19908 = w19833 ^ w19807;
	assign w19797 = w19855 ^ w19828;
	assign w49041 = w19796 ^ w19797;
	assign w19810 = w19814 ^ w44200;
	assign w19809 = w19805 ^ w19810;
	assign w19909 = w19808 ^ w19809;
	assign w44203 = w19853 ^ w19854;
	assign w49042 = w44203 ^ w19833;
	assign w19835 = w19850 ^ w44203;
	assign w19801 = w19846 ^ w19835;
	assign w19798 = ~w19801;
	assign w19795 = w19851 ^ w19835;
	assign w49043 = w19824 ^ w19795;
	assign w44204 = w19855 ^ w19857;
	assign w19813 = w44204 ^ w19810;
	assign w19910 = w19812 ^ w19813;
	assign w19800 = w19804 ^ w44204;
	assign w19803 = w19842 ^ w19800;
	assign w19907 = w19802 ^ w19803;
	assign w19799 = w19823 ^ w19800;
	assign w49040 = w19798 ^ w19799;
	assign w44688 = w31539 ^ w31545;
	assign w31451 = w31483 ^ w44688;
	assign w31494 = w47447 ^ w31451;
	assign w31529 = w31534 ^ w31494;
	assign w31489 = w44688 ^ w31474;
	assign w31535 = w31497 ^ w31489;
	assign w44689 = w31539 ^ w31542;
	assign w31492 = w31540 ^ w44689;
	assign w31448 = w31543 ^ w31492;
	assign w31530 = w47451 ^ w31448;
	assign w31528 = w31529 & w31530;
	assign w31446 = w31528 ^ w31545;
	assign w31526 = w31534 ^ w31528;
	assign w31441 = w31446 ^ w31542;
	assign w31447 = w31528 ^ w31492;
	assign w31452 = w31478 ^ w44689;
	assign w31536 = w31452 ^ w31477;
	assign w31527 = w31528 ^ w31536;
	assign w31533 = w31534 ^ w31536;
	assign w31532 = w31535 & w31533;
	assign w31531 = w31532 ^ w31494;
	assign w31443 = w31532 ^ w31544;
	assign w31439 = w31443 ^ w31479;
	assign w31442 = w47445 ^ w31439;
	assign w31519 = w31441 ^ w31442;
	assign w31440 = w31532 ^ w31488;
	assign w31438 = w47447 ^ w31439;
	assign w31525 = w31536 & w31526;
	assign w31523 = w31525 ^ w31533;
	assign w31522 = w31531 & w31523;
	assign w31487 = w31522 ^ w31497;
	assign w31521 = w31487 ^ w31489;
	assign w31445 = w31522 ^ w31546;
	assign w31518 = w31487 ^ w31440;
	assign w31513 = w31527 & w47452;
	assign w31512 = w31518 & w31548;
	assign w31511 = w31521 & w31560;
	assign w31510 = w31531 & w31550;
	assign w31454 = w31510 ^ w31511;
	assign w31509 = w31519 & w31551;
	assign w31504 = w31527 & w31559;
	assign w31503 = w31518 & w31563;
	assign w31470 = w31512 ^ w31503;
	assign w31502 = w31521 & w31556;
	assign w31472 = w31510 ^ w31502;
	assign w31501 = w31531 & w31557;
	assign w31500 = w31519 & w31562;
	assign w44691 = w31511 ^ w31512;
	assign w44693 = w31525 ^ w31543;
	assign w31517 = w44693 ^ w31495;
	assign w31515 = w31517 & w31554;
	assign w44692 = w31513 ^ w31515;
	assign w31506 = w31517 & w31558;
	assign w31484 = w47451 ^ w44693;
	assign w31524 = w31484 ^ w31447;
	assign w31437 = w31484 ^ w31445;
	assign w31444 = w31474 ^ w31437;
	assign w31520 = w31441 ^ w31444;
	assign w31516 = w31437 ^ w31438;
	assign w31514 = w31524 & w31553;
	assign w31508 = w31516 & w31549;
	assign w31493 = w31508 ^ w44691;
	assign w31469 = w31508 ^ w31511;
	assign w31466 = ~w31469;
	assign w31465 = w31508 ^ w31509;
	assign w31459 = w31504 ^ w31493;
	assign w31456 = ~w31459;
	assign w31453 = w31509 ^ w31493;
	assign w31507 = w31520 & w31552;
	assign w31485 = w31503 ^ w31507;
	assign w31463 = ~w31485;
	assign w31462 = w31463 ^ w31501;
	assign w31458 = w31462 ^ w44692;
	assign w31461 = w31500 ^ w31458;
	assign w31505 = w31524 & w31555;
	assign w31499 = w31516 & w31564;
	assign w31498 = w31520 & w31561;
	assign w31464 = w31509 ^ w31498;
	assign w31460 = ~w31464;
	assign w31565 = w31460 ^ w31461;
	assign w44690 = w31499 ^ w31500;
	assign w31481 = w31505 ^ w44690;
	assign w31457 = w31481 ^ w31458;
	assign w49073 = w31456 ^ w31457;
	assign w31482 = w31506 ^ w31481;
	assign w49076 = w31482 ^ w31453;
	assign w31486 = w31514 ^ w31482;
	assign w31455 = w31513 ^ w31486;
	assign w49074 = w31454 ^ w31455;
	assign w31491 = w31515 ^ w31486;
	assign w31566 = w31491 ^ w31465;
	assign w7501 = w49063 ^ w49076;
	assign w7252 = w7501 ^ w49074;
	assign w7248 = ~w7501;
	assign w7249 = w7248 ^ w49073;
	assign w49075 = w44691 ^ w31491;
	assign w31468 = w31472 ^ w44690;
	assign w31471 = w44692 ^ w31468;
	assign w31568 = w31470 ^ w31471;
	assign w31467 = w31463 ^ w31468;
	assign w31567 = w31466 ^ w31467;
	assign w6915 = w45465 ^ w45273;
	assign w7231 = w6914 ^ w6915;
	assign w48760 = w7231 ^ w7187;
	assign w47459 = w48760 ^ w1422;
	assign w19681 = w47459 ^ w47457;
	assign w19683 = w47458 ^ w19681;
	assign w19759 = w47454 ^ w19683;
	assign w19756 = w47455 ^ w19683;
	assign w19758 = w19688 ^ w19683;
	assign w19764 = w47459 ^ w19768;
	assign w19762 = w19681 ^ w19770;
	assign w19761 = w47460 ^ w19762;
	assign w19698 = w47459 ^ w47458;
	assign w19763 = w19698 ^ w19765;
	assign w19766 = w19770 ^ w19698;
	assign w19760 = w19681 ^ w19644;
	assign w19771 = w47453 ^ w47459;
	assign w19755 = w19762 & w19766;
	assign w19687 = w19755 ^ w19684;
	assign w19754 = w19763 & w19761;
	assign w19705 = w19748 ^ w19754;
	assign w19752 = w19771 & w19756;
	assign w19686 = w19752 ^ w19682;
	assign w19751 = w19768 & w19764;
	assign w19750 = w19765 & w19758;
	assign w19749 = w19770 & w19759;
	assign w19685 = w19749 ^ w19683;
	assign w19691 = w19687 ^ w19685;
	assign w19696 = w47453 ^ w19691;
	assign w19746 = w19705 ^ w19696;
	assign w19657 = w19748 ^ w19749;
	assign w19704 = w19657 ^ w19658;
	assign w19703 = w19704 ^ w19686;
	assign w19745 = w19751 ^ w19703;
	assign w19747 = w19769 & w19760;
	assign w19742 = w19746 & w19745;
	assign w44193 = w19747 ^ w19753;
	assign w19659 = w19691 ^ w44193;
	assign w19702 = w47455 ^ w19659;
	assign w19737 = w19742 ^ w19702;
	assign w19697 = w44193 ^ w19682;
	assign w19743 = w19705 ^ w19697;
	assign w44194 = w19747 ^ w19750;
	assign w19700 = w19748 ^ w44194;
	assign w19656 = w19751 ^ w19700;
	assign w19738 = w47459 ^ w19656;
	assign w19736 = w19737 & w19738;
	assign w19655 = w19736 ^ w19700;
	assign w19734 = w19742 ^ w19736;
	assign w19654 = w19736 ^ w19753;
	assign w19649 = w19654 ^ w19750;
	assign w19660 = w19686 ^ w44194;
	assign w19744 = w19660 ^ w19685;
	assign w19735 = w19736 ^ w19744;
	assign w19741 = w19742 ^ w19744;
	assign w19740 = w19743 & w19741;
	assign w19739 = w19740 ^ w19702;
	assign w19651 = w19740 ^ w19752;
	assign w19647 = w19651 ^ w19687;
	assign w19650 = w47453 ^ w19647;
	assign w19727 = w19649 ^ w19650;
	assign w19648 = w19740 ^ w19696;
	assign w19646 = w47455 ^ w19647;
	assign w19733 = w19744 & w19734;
	assign w19731 = w19733 ^ w19741;
	assign w19730 = w19739 & w19731;
	assign w19695 = w19730 ^ w19705;
	assign w19729 = w19695 ^ w19697;
	assign w19653 = w19730 ^ w19754;
	assign w19726 = w19695 ^ w19648;
	assign w19721 = w19735 & w47460;
	assign w19720 = w19726 & w19756;
	assign w19719 = w19729 & w19768;
	assign w19718 = w19739 & w19758;
	assign w19662 = w19718 ^ w19719;
	assign w19717 = w19727 & w19759;
	assign w19712 = w19735 & w19767;
	assign w19711 = w19726 & w19771;
	assign w19678 = w19720 ^ w19711;
	assign w19710 = w19729 & w19764;
	assign w19680 = w19718 ^ w19710;
	assign w19709 = w19739 & w19765;
	assign w19708 = w19727 & w19770;
	assign w44196 = w19719 ^ w19720;
	assign w44198 = w19733 ^ w19751;
	assign w19725 = w44198 ^ w19703;
	assign w19723 = w19725 & w19762;
	assign w44197 = w19721 ^ w19723;
	assign w19714 = w19725 & w19766;
	assign w19692 = w47459 ^ w44198;
	assign w19732 = w19692 ^ w19655;
	assign w19645 = w19692 ^ w19653;
	assign w19652 = w19682 ^ w19645;
	assign w19728 = w19649 ^ w19652;
	assign w19724 = w19645 ^ w19646;
	assign w19722 = w19732 & w19761;
	assign w19716 = w19724 & w19757;
	assign w19701 = w19716 ^ w44196;
	assign w19677 = w19716 ^ w19719;
	assign w19674 = ~w19677;
	assign w19673 = w19716 ^ w19717;
	assign w19667 = w19712 ^ w19701;
	assign w19664 = ~w19667;
	assign w19661 = w19717 ^ w19701;
	assign w19715 = w19728 & w19760;
	assign w19693 = w19711 ^ w19715;
	assign w19671 = ~w19693;
	assign w19670 = w19671 ^ w19709;
	assign w19666 = w19670 ^ w44197;
	assign w19669 = w19708 ^ w19666;
	assign w19713 = w19732 & w19763;
	assign w19707 = w19724 & w19772;
	assign w19706 = w19728 & w19769;
	assign w19672 = w19717 ^ w19706;
	assign w19668 = ~w19672;
	assign w19773 = w19668 ^ w19669;
	assign w44195 = w19707 ^ w19708;
	assign w19689 = w19713 ^ w44195;
	assign w19665 = w19689 ^ w19666;
	assign w49088 = w19664 ^ w19665;
	assign w19690 = w19714 ^ w19689;
	assign w49091 = w19690 ^ w19661;
	assign w19694 = w19722 ^ w19690;
	assign w19663 = w19721 ^ w19694;
	assign w49089 = w19662 ^ w19663;
	assign w19699 = w19723 ^ w19694;
	assign w19774 = w19699 ^ w19673;
	assign w49090 = w44196 ^ w19699;
	assign w19676 = w19680 ^ w44195;
	assign w19679 = w44197 ^ w19676;
	assign w19776 = w19678 ^ w19679;
	assign w19675 = w19671 ^ w19676;
	assign w19775 = w19674 ^ w19675;
	assign w45434 = ~w19775;
	assign w45435 = ~w19776;
	assign w45438 = ~w19909;
	assign w45439 = ~w19910;
	assign w45440 = ~w19773;
	assign w45441 = ~w19774;
	assign w45444 = ~w19907;
	assign w45445 = ~w19908;
	assign w45546 = ~w25134;
	assign w7383 = w49063 ^ w45546;
	assign w45547 = ~w25135;
	assign w45548 = ~w25136;
	assign w45553 = ~w25133;
	assign w45726 = ~w31566;
	assign w7510 = w45546 ^ w45726;
	assign w45727 = ~w31567;
	assign w45728 = ~w31568;
	assign w7246 = w7248 ^ w45728;
	assign w45733 = ~w31565;
	assign w7402 = w45733 ^ w45553;
	assign w45887 = ~w7149;
	assign w6971 = w45887 ^ w48894;
	assign w48798 = w6971 ^ w6972;
	assign w6994 = w45887 ^ w45194;
	assign w6990 = w45887 ^ w48877;
	assign w48786 = w6989 ^ w6990;
	assign w6992 = w6993 ^ w6994;
	assign w48784 = ~w6992;
	assign w47421 = w48798 ^ w1396;
	assign w19548 = w47423 ^ w47421;
	assign w19623 = w19548 ^ w19638;
	assign w19636 = w47424 ^ w47421;
	assign w19632 = w19636 ^ w19564;
	assign w19631 = w19548 ^ w19554;
	assign w19629 = w19564 ^ w19631;
	assign w19628 = w19547 ^ w19636;
	assign w19627 = w47428 ^ w19628;
	assign w19510 = w19550 ^ w19548;
	assign w19626 = w19547 ^ w19510;
	assign w19637 = w47421 ^ w47427;
	assign w19635 = w47421 ^ w47426;
	assign w19621 = w19628 & w19632;
	assign w19553 = w19621 ^ w19550;
	assign w19620 = w19629 & w19627;
	assign w19618 = w19637 & w19622;
	assign w19552 = w19618 ^ w19548;
	assign w19616 = w19631 & w19624;
	assign w19615 = w19636 & w19625;
	assign w19551 = w19615 ^ w19549;
	assign w19557 = w19553 ^ w19551;
	assign w19562 = w47421 ^ w19557;
	assign w19614 = w19638 & w19623;
	assign w19571 = w19614 ^ w19620;
	assign w19612 = w19571 ^ w19562;
	assign w19523 = w19614 ^ w19615;
	assign w19570 = w19523 ^ w19524;
	assign w19569 = w19570 ^ w19552;
	assign w19611 = w19617 ^ w19569;
	assign w19613 = w19635 & w19626;
	assign w19608 = w19612 & w19611;
	assign w47435 = w48784 ^ w1382;
	assign w13473 = w47429 ^ w47435;
	assign w13466 = w47435 ^ w13470;
	assign w47433 = w48786 ^ w1384;
	assign w13360 = w47433 ^ w47434;
	assign w13383 = w47435 ^ w47433;
	assign w13385 = w47434 ^ w13383;
	assign w13460 = w13390 ^ w13385;
	assign w13452 = w13467 & w13460;
	assign w13461 = w47430 ^ w13385;
	assign w6988 = w45887 ^ w48878;
	assign w48787 = w6987 ^ w6988;
	assign w47432 = w48787 ^ w1385;
	assign w13474 = w47434 ^ w47432;
	assign w13459 = w13384 ^ w13474;
	assign w13450 = w13474 & w13459;
	assign w13386 = w47432 ^ w47430;
	assign w13346 = w13386 ^ w13384;
	assign w13345 = w13386 ^ w47431;
	assign w13462 = w13383 ^ w13346;
	assign w13469 = w47436 ^ w13345;
	assign w13455 = w47436 & w13469;
	assign w13472 = w47432 ^ w47429;
	assign w13451 = w13472 & w13461;
	assign w13359 = w13450 ^ w13451;
	assign w13406 = w13359 ^ w13360;
	assign w13387 = w13451 ^ w13385;
	assign w13464 = w13383 ^ w13472;
	assign w13463 = w47436 ^ w13464;
	assign w13458 = w47431 ^ w13385;
	assign w13454 = w13473 & w13458;
	assign w13388 = w13454 ^ w13384;
	assign w13405 = w13406 ^ w13388;
	assign w13453 = w13470 & w13466;
	assign w13447 = w13453 ^ w13405;
	assign w44188 = w19613 ^ w19619;
	assign w19563 = w44188 ^ w19548;
	assign w19609 = w19571 ^ w19563;
	assign w19525 = w19557 ^ w44188;
	assign w19568 = w47423 ^ w19525;
	assign w19603 = w19608 ^ w19568;
	assign w44189 = w19613 ^ w19616;
	assign w19566 = w19614 ^ w44189;
	assign w19522 = w19617 ^ w19566;
	assign w19604 = w47427 ^ w19522;
	assign w19602 = w19603 & w19604;
	assign w19521 = w19602 ^ w19566;
	assign w19520 = w19602 ^ w19619;
	assign w19515 = w19520 ^ w19616;
	assign w19600 = w19608 ^ w19602;
	assign w19526 = w19552 ^ w44189;
	assign w19610 = w19526 ^ w19551;
	assign w19601 = w19602 ^ w19610;
	assign w19607 = w19608 ^ w19610;
	assign w19606 = w19609 & w19607;
	assign w19605 = w19606 ^ w19568;
	assign w19517 = w19606 ^ w19618;
	assign w19513 = w19517 ^ w19553;
	assign w19516 = w47421 ^ w19513;
	assign w19593 = w19515 ^ w19516;
	assign w19514 = w19606 ^ w19562;
	assign w19512 = w47423 ^ w19513;
	assign w19599 = w19610 & w19600;
	assign w19597 = w19599 ^ w19607;
	assign w19596 = w19605 & w19597;
	assign w19561 = w19596 ^ w19571;
	assign w19595 = w19561 ^ w19563;
	assign w19519 = w19596 ^ w19620;
	assign w19592 = w19561 ^ w19514;
	assign w19587 = w19601 & w47428;
	assign w19586 = w19592 & w19622;
	assign w19585 = w19595 & w19634;
	assign w19584 = w19605 & w19624;
	assign w19528 = w19584 ^ w19585;
	assign w19583 = w19593 & w19625;
	assign w19578 = w19601 & w19633;
	assign w19577 = w19592 & w19637;
	assign w19544 = w19586 ^ w19577;
	assign w19576 = w19595 & w19630;
	assign w19546 = w19584 ^ w19576;
	assign w19575 = w19605 & w19631;
	assign w19574 = w19593 & w19636;
	assign w44190 = w19585 ^ w19586;
	assign w44192 = w19599 ^ w19617;
	assign w19558 = w47427 ^ w44192;
	assign w19598 = w19558 ^ w19521;
	assign w19579 = w19598 & w19629;
	assign w19588 = w19598 & w19627;
	assign w19511 = w19558 ^ w19519;
	assign w19518 = w19548 ^ w19511;
	assign w19594 = w19515 ^ w19518;
	assign w19581 = w19594 & w19626;
	assign w19559 = w19577 ^ w19581;
	assign w19537 = ~w19559;
	assign w19536 = w19537 ^ w19575;
	assign w19590 = w19511 ^ w19512;
	assign w19573 = w19590 & w19638;
	assign w19572 = w19594 & w19635;
	assign w19538 = w19583 ^ w19572;
	assign w19534 = ~w19538;
	assign w43553 = w19573 ^ w19574;
	assign w19555 = w19579 ^ w43553;
	assign w19542 = w19546 ^ w43553;
	assign w19541 = w19537 ^ w19542;
	assign w19582 = w19590 & w19623;
	assign w19539 = w19582 ^ w19583;
	assign w19567 = w19582 ^ w44190;
	assign w19533 = w19578 ^ w19567;
	assign w19530 = ~w19533;
	assign w19527 = w19583 ^ w19567;
	assign w19543 = w19582 ^ w19585;
	assign w19540 = ~w19543;
	assign w19641 = w19540 ^ w19541;
	assign w19591 = w44192 ^ w19569;
	assign w19589 = w19591 & w19628;
	assign w19580 = w19591 & w19632;
	assign w19556 = w19580 ^ w19555;
	assign w19560 = w19588 ^ w19556;
	assign w19565 = w19589 ^ w19560;
	assign w49107 = w44190 ^ w19565;
	assign w19640 = w19565 ^ w19539;
	assign w19529 = w19587 ^ w19560;
	assign w49106 = w19528 ^ w19529;
	assign w49108 = w19556 ^ w19527;
	assign w7296 = w49107 ^ w49106;
	assign w44191 = w19587 ^ w19589;
	assign w19545 = w44191 ^ w19542;
	assign w19642 = w19544 ^ w19545;
	assign w19532 = w19536 ^ w44191;
	assign w19535 = w19574 ^ w19532;
	assign w19639 = w19534 ^ w19535;
	assign w19531 = w19555 ^ w19532;
	assign w49105 = w19530 ^ w19531;
	assign w13400 = w47435 ^ w47434;
	assign w13465 = w13400 ^ w13467;
	assign w13456 = w13465 & w13463;
	assign w13468 = w13472 ^ w13400;
	assign w13457 = w13464 & w13468;
	assign w13389 = w13457 ^ w13386;
	assign w13393 = w13389 ^ w13387;
	assign w13407 = w13450 ^ w13456;
	assign w13398 = w47429 ^ w13393;
	assign w13448 = w13407 ^ w13398;
	assign w13449 = w13471 & w13462;
	assign w43931 = w13449 ^ w13452;
	assign w13362 = w13388 ^ w43931;
	assign w13446 = w13362 ^ w13387;
	assign w13402 = w13450 ^ w43931;
	assign w13358 = w13453 ^ w13402;
	assign w13440 = w47435 ^ w13358;
	assign w43934 = w13449 ^ w13455;
	assign w13361 = w13393 ^ w43934;
	assign w13404 = w47431 ^ w13361;
	assign w13399 = w43934 ^ w13384;
	assign w13445 = w13407 ^ w13399;
	assign w13444 = w13448 & w13447;
	assign w13443 = w13444 ^ w13446;
	assign w13442 = w13445 & w13443;
	assign w13350 = w13442 ^ w13398;
	assign w13353 = w13442 ^ w13454;
	assign w13349 = w13353 ^ w13389;
	assign w13348 = w47431 ^ w13349;
	assign w13352 = w47429 ^ w13349;
	assign w13439 = w13444 ^ w13404;
	assign w13438 = w13439 & w13440;
	assign w13356 = w13438 ^ w13455;
	assign w13351 = w13356 ^ w13452;
	assign w13357 = w13438 ^ w13402;
	assign w13429 = w13351 ^ w13352;
	assign w13419 = w13429 & w13461;
	assign w13436 = w13444 ^ w13438;
	assign w13435 = w13446 & w13436;
	assign w13441 = w13442 ^ w13404;
	assign w13420 = w13441 & w13460;
	assign w13411 = w13441 & w13467;
	assign w13433 = w13435 ^ w13443;
	assign w13432 = w13441 & w13433;
	assign w13355 = w13432 ^ w13456;
	assign w13410 = w13429 & w13472;
	assign w13437 = w13438 ^ w13446;
	assign w13423 = w13437 & w47436;
	assign w13414 = w13437 & w13469;
	assign w13397 = w13432 ^ w13407;
	assign w13428 = w13397 ^ w13350;
	assign w13422 = w13428 & w13458;
	assign w13431 = w13397 ^ w13399;
	assign w13421 = w13431 & w13470;
	assign w13364 = w13420 ^ w13421;
	assign w13413 = w13428 & w13473;
	assign w13380 = w13422 ^ w13413;
	assign w13412 = w13431 & w13466;
	assign w43933 = w13435 ^ w13453;
	assign w13427 = w43933 ^ w13405;
	assign w13416 = w13427 & w13468;
	assign w13425 = w13427 & w13464;
	assign w13394 = w47435 ^ w43933;
	assign w13434 = w13394 ^ w13357;
	assign w13347 = w13394 ^ w13355;
	assign w13354 = w13384 ^ w13347;
	assign w13424 = w13434 & w13463;
	assign w13430 = w13351 ^ w13354;
	assign w13408 = w13430 & w13471;
	assign w13417 = w13430 & w13462;
	assign w13374 = w13419 ^ w13408;
	assign w13370 = ~w13374;
	assign w13426 = w13347 ^ w13348;
	assign w13418 = w13426 & w13459;
	assign w13379 = w13418 ^ w13421;
	assign w13375 = w13418 ^ w13419;
	assign w13376 = ~w13379;
	assign w13395 = w13413 ^ w13417;
	assign w13373 = ~w13395;
	assign w13372 = w13373 ^ w13411;
	assign w13415 = w13434 & w13465;
	assign w43935 = w13421 ^ w13422;
	assign w13403 = w13418 ^ w43935;
	assign w13369 = w13414 ^ w13403;
	assign w13363 = w13419 ^ w13403;
	assign w13366 = ~w13369;
	assign w43936 = w13423 ^ w13425;
	assign w13368 = w13372 ^ w43936;
	assign w13371 = w13410 ^ w13368;
	assign w13475 = w13370 ^ w13371;
	assign w49047 = ~w13475;
	assign w7547 = w45444 ^ w49047;
	assign w13382 = w13420 ^ w13412;
	assign w13409 = w13426 & w13474;
	assign w43932 = w13409 ^ w13410;
	assign w13391 = w13415 ^ w43932;
	assign w13392 = w13416 ^ w13391;
	assign w49049 = w13392 ^ w13363;
	assign w13396 = w13424 ^ w13392;
	assign w13401 = w13425 ^ w13396;
	assign w13365 = w13423 ^ w13396;
	assign w49045 = w13364 ^ w13365;
	assign w13476 = w13401 ^ w13375;
	assign w49048 = ~w13476;
	assign w49046 = w43935 ^ w13401;
	assign w7495 = w49043 ^ w49049;
	assign w7285 = w7495 ^ w49041;
	assign w7550 = w49042 ^ w49046;
	assign w7559 = w49041 ^ w49045;
	assign w7545 = w45445 ^ w49048;
	assign w7441 = ~w7559;
	assign w13367 = w13391 ^ w13368;
	assign w49044 = w13366 ^ w13367;
	assign w7286 = w49040 ^ w49044;
	assign w7564 = w7285 ^ w7286;
	assign w13378 = w13382 ^ w43932;
	assign w13381 = w43936 ^ w13378;
	assign w13478 = w13380 ^ w13381;
	assign w13377 = w13373 ^ w13378;
	assign w13477 = w13376 ^ w13377;
	assign w45267 = ~w13477;
	assign w45268 = ~w13478;
	assign w45430 = ~w19641;
	assign w45431 = ~w19642;
	assign w45436 = ~w19639;
	assign w45437 = ~w19640;
	assign w7444 = w45437 ^ w45436;
	assign w45908 = ~w6671;
	assign w6466 = w45908 ^ w48653;
	assign w6739 = w6466 ^ w6467;
	assign w48537 = w6739 ^ w6736;
	assign w47609 = w48537 ^ w2005;
	assign w28659 = w47611 ^ w47609;
	assign w28661 = w47610 ^ w28659;
	assign w28737 = w47606 ^ w28661;
	assign w28734 = w47607 ^ w28661;
	assign w28736 = w28666 ^ w28661;
	assign w28636 = w47609 ^ w47610;
	assign w28730 = w28749 & w28734;
	assign w28664 = w28730 ^ w28660;
	assign w28728 = w28743 & w28736;
	assign w6503 = w45908 ^ w45656;
	assign w48517 = w6503 ^ w6504;
	assign w47629 = w48517 ^ w1985;
	assign w25444 = w47631 ^ w47629;
	assign w25519 = w25444 ^ w25534;
	assign w25532 = w47632 ^ w47629;
	assign w25528 = w25532 ^ w25460;
	assign w25527 = w25444 ^ w25450;
	assign w25525 = w25460 ^ w25527;
	assign w25524 = w25443 ^ w25532;
	assign w25523 = w47636 ^ w25524;
	assign w25406 = w25446 ^ w25444;
	assign w25522 = w25443 ^ w25406;
	assign w25533 = w47629 ^ w47635;
	assign w25531 = w47629 ^ w47634;
	assign w25517 = w25524 & w25528;
	assign w25449 = w25517 ^ w25446;
	assign w25516 = w25525 & w25523;
	assign w25514 = w25533 & w25518;
	assign w25448 = w25514 ^ w25444;
	assign w25512 = w25527 & w25520;
	assign w25511 = w25532 & w25521;
	assign w25447 = w25511 ^ w25445;
	assign w25453 = w25449 ^ w25447;
	assign w25458 = w47629 ^ w25453;
	assign w25510 = w25534 & w25519;
	assign w25467 = w25510 ^ w25516;
	assign w25508 = w25467 ^ w25458;
	assign w25419 = w25510 ^ w25511;
	assign w25466 = w25419 ^ w25420;
	assign w25465 = w25466 ^ w25448;
	assign w25507 = w25513 ^ w25465;
	assign w25509 = w25531 & w25522;
	assign w25504 = w25508 & w25507;
	assign w6590 = w45908 ^ w48651;
	assign w48538 = w6589 ^ w6590;
	assign w47608 = w48538 ^ w2006;
	assign w28662 = w47608 ^ w47606;
	assign w28748 = w47608 ^ w47605;
	assign w28744 = w28748 ^ w28676;
	assign w28740 = w28659 ^ w28748;
	assign w28739 = w47612 ^ w28740;
	assign w28750 = w47610 ^ w47608;
	assign w28735 = w28660 ^ w28750;
	assign w28622 = w28662 ^ w28660;
	assign w28738 = w28659 ^ w28622;
	assign w28621 = w28662 ^ w47607;
	assign w28745 = w47612 ^ w28621;
	assign w28733 = w28740 & w28744;
	assign w28665 = w28733 ^ w28662;
	assign w28732 = w28741 & w28739;
	assign w28731 = w47612 & w28745;
	assign w28727 = w28748 & w28737;
	assign w28663 = w28727 ^ w28661;
	assign w28669 = w28665 ^ w28663;
	assign w28674 = w47605 ^ w28669;
	assign w28726 = w28750 & w28735;
	assign w28683 = w28726 ^ w28732;
	assign w28724 = w28683 ^ w28674;
	assign w28635 = w28726 ^ w28727;
	assign w28682 = w28635 ^ w28636;
	assign w28681 = w28682 ^ w28664;
	assign w28723 = w28729 ^ w28681;
	assign w28725 = w28747 & w28738;
	assign w28720 = w28724 & w28723;
	assign w44435 = w25509 ^ w25515;
	assign w25459 = w44435 ^ w25444;
	assign w25505 = w25467 ^ w25459;
	assign w25421 = w25453 ^ w44435;
	assign w25464 = w47631 ^ w25421;
	assign w25499 = w25504 ^ w25464;
	assign w44436 = w25509 ^ w25512;
	assign w25462 = w25510 ^ w44436;
	assign w25418 = w25513 ^ w25462;
	assign w25500 = w47635 ^ w25418;
	assign w25498 = w25499 & w25500;
	assign w25496 = w25504 ^ w25498;
	assign w25417 = w25498 ^ w25462;
	assign w25416 = w25498 ^ w25515;
	assign w25411 = w25416 ^ w25512;
	assign w25422 = w25448 ^ w44436;
	assign w25506 = w25422 ^ w25447;
	assign w25497 = w25498 ^ w25506;
	assign w25503 = w25504 ^ w25506;
	assign w25502 = w25505 & w25503;
	assign w25501 = w25502 ^ w25464;
	assign w25413 = w25502 ^ w25514;
	assign w25409 = w25413 ^ w25449;
	assign w25412 = w47629 ^ w25409;
	assign w25489 = w25411 ^ w25412;
	assign w25410 = w25502 ^ w25458;
	assign w25408 = w47631 ^ w25409;
	assign w25495 = w25506 & w25496;
	assign w25493 = w25495 ^ w25503;
	assign w25492 = w25501 & w25493;
	assign w25457 = w25492 ^ w25467;
	assign w25491 = w25457 ^ w25459;
	assign w25415 = w25492 ^ w25516;
	assign w25488 = w25457 ^ w25410;
	assign w25483 = w25497 & w47636;
	assign w25482 = w25488 & w25518;
	assign w25481 = w25491 & w25530;
	assign w25480 = w25501 & w25520;
	assign w25424 = w25480 ^ w25481;
	assign w25479 = w25489 & w25521;
	assign w25474 = w25497 & w25529;
	assign w25473 = w25488 & w25533;
	assign w25440 = w25482 ^ w25473;
	assign w25472 = w25491 & w25526;
	assign w25442 = w25480 ^ w25472;
	assign w25471 = w25501 & w25527;
	assign w25470 = w25489 & w25532;
	assign w44437 = w25481 ^ w25482;
	assign w44439 = w25495 ^ w25513;
	assign w25454 = w47635 ^ w44439;
	assign w25407 = w25454 ^ w25415;
	assign w25414 = w25444 ^ w25407;
	assign w25490 = w25411 ^ w25414;
	assign w25477 = w25490 & w25522;
	assign w25455 = w25473 ^ w25477;
	assign w25433 = ~w25455;
	assign w25486 = w25407 ^ w25408;
	assign w25478 = w25486 & w25519;
	assign w25435 = w25478 ^ w25479;
	assign w25439 = w25478 ^ w25481;
	assign w25436 = ~w25439;
	assign w25432 = w25433 ^ w25471;
	assign w25469 = w25486 & w25534;
	assign w25468 = w25490 & w25531;
	assign w25434 = w25479 ^ w25468;
	assign w25430 = ~w25434;
	assign w43570 = w25469 ^ w25470;
	assign w25438 = w25442 ^ w43570;
	assign w25437 = w25433 ^ w25438;
	assign w25537 = w25436 ^ w25437;
	assign w25494 = w25454 ^ w25417;
	assign w25484 = w25494 & w25523;
	assign w25475 = w25494 & w25525;
	assign w25451 = w25475 ^ w43570;
	assign w25463 = w25478 ^ w44437;
	assign w25429 = w25474 ^ w25463;
	assign w25426 = ~w25429;
	assign w25423 = w25479 ^ w25463;
	assign w25487 = w44439 ^ w25465;
	assign w25485 = w25487 & w25524;
	assign w25476 = w25487 & w25528;
	assign w25452 = w25476 ^ w25451;
	assign w25456 = w25484 ^ w25452;
	assign w25461 = w25485 ^ w25456;
	assign w48897 = w44437 ^ w25461;
	assign w25536 = w25461 ^ w25435;
	assign w25425 = w25483 ^ w25456;
	assign w48896 = w25424 ^ w25425;
	assign w48899 = w25452 ^ w25423;
	assign w48898 = ~w25536;
	assign w7156 = w48899 ^ w48911;
	assign w6955 = w7194 ^ w7156;
	assign w7170 = w48896 ^ w48909;
	assign w6950 = ~w48897;
	assign w7139 = w48910 ^ w6950;
	assign w44438 = w25483 ^ w25485;
	assign w25441 = w44438 ^ w25438;
	assign w25538 = w25440 ^ w25441;
	assign w25428 = w25432 ^ w44438;
	assign w25431 = w25470 ^ w25428;
	assign w25535 = w25430 ^ w25431;
	assign w25427 = w25451 ^ w25428;
	assign w48895 = w25426 ^ w25427;
	assign w6912 = w7156 ^ w48895;
	assign w7232 = w6912 ^ w6913;
	assign w44569 = w28725 ^ w28731;
	assign w28675 = w44569 ^ w28660;
	assign w28721 = w28683 ^ w28675;
	assign w28637 = w28669 ^ w44569;
	assign w28680 = w47607 ^ w28637;
	assign w28715 = w28720 ^ w28680;
	assign w44570 = w28725 ^ w28728;
	assign w28678 = w28726 ^ w44570;
	assign w28634 = w28729 ^ w28678;
	assign w28716 = w47611 ^ w28634;
	assign w28714 = w28715 & w28716;
	assign w28633 = w28714 ^ w28678;
	assign w28632 = w28714 ^ w28731;
	assign w28627 = w28632 ^ w28728;
	assign w28712 = w28720 ^ w28714;
	assign w28638 = w28664 ^ w44570;
	assign w28722 = w28638 ^ w28663;
	assign w28713 = w28714 ^ w28722;
	assign w28719 = w28720 ^ w28722;
	assign w28718 = w28721 & w28719;
	assign w28717 = w28718 ^ w28680;
	assign w28629 = w28718 ^ w28730;
	assign w28625 = w28629 ^ w28665;
	assign w28628 = w47605 ^ w28625;
	assign w28705 = w28627 ^ w28628;
	assign w28626 = w28718 ^ w28674;
	assign w28624 = w47607 ^ w28625;
	assign w28711 = w28722 & w28712;
	assign w28709 = w28711 ^ w28719;
	assign w28708 = w28717 & w28709;
	assign w28673 = w28708 ^ w28683;
	assign w28707 = w28673 ^ w28675;
	assign w28631 = w28708 ^ w28732;
	assign w28704 = w28673 ^ w28626;
	assign w28699 = w28713 & w47612;
	assign w28698 = w28704 & w28734;
	assign w28697 = w28707 & w28746;
	assign w28696 = w28717 & w28736;
	assign w28640 = w28696 ^ w28697;
	assign w28695 = w28705 & w28737;
	assign w28690 = w28713 & w28745;
	assign w28689 = w28704 & w28749;
	assign w28656 = w28698 ^ w28689;
	assign w28688 = w28707 & w28742;
	assign w28658 = w28696 ^ w28688;
	assign w28687 = w28717 & w28743;
	assign w28686 = w28705 & w28748;
	assign w44571 = w28697 ^ w28698;
	assign w44573 = w28711 ^ w28729;
	assign w28670 = w47611 ^ w44573;
	assign w28710 = w28670 ^ w28633;
	assign w28691 = w28710 & w28741;
	assign w28700 = w28710 & w28739;
	assign w28623 = w28670 ^ w28631;
	assign w28630 = w28660 ^ w28623;
	assign w28706 = w28627 ^ w28630;
	assign w28693 = w28706 & w28738;
	assign w28671 = w28689 ^ w28693;
	assign w28649 = ~w28671;
	assign w28648 = w28649 ^ w28687;
	assign w28702 = w28623 ^ w28624;
	assign w28685 = w28702 & w28750;
	assign w28684 = w28706 & w28747;
	assign w28650 = w28695 ^ w28684;
	assign w28646 = ~w28650;
	assign w43580 = w28685 ^ w28686;
	assign w28654 = w28658 ^ w43580;
	assign w28653 = w28649 ^ w28654;
	assign w28667 = w28691 ^ w43580;
	assign w28694 = w28702 & w28735;
	assign w28651 = w28694 ^ w28695;
	assign w28679 = w28694 ^ w44571;
	assign w28645 = w28690 ^ w28679;
	assign w28642 = ~w28645;
	assign w28639 = w28695 ^ w28679;
	assign w28655 = w28694 ^ w28697;
	assign w28652 = ~w28655;
	assign w28753 = w28652 ^ w28653;
	assign w28703 = w44573 ^ w28681;
	assign w28701 = w28703 & w28740;
	assign w28692 = w28703 & w28744;
	assign w28668 = w28692 ^ w28667;
	assign w28672 = w28700 ^ w28668;
	assign w28677 = w28701 ^ w28672;
	assign w48856 = w44571 ^ w28677;
	assign w28752 = w28677 ^ w28651;
	assign w28641 = w28699 ^ w28672;
	assign w48855 = w28640 ^ w28641;
	assign w7085 = w7086 ^ w48855;
	assign w48858 = w28668 ^ w28639;
	assign w48857 = ~w28752;
	assign w48730 = w7084 ^ w7085;
	assign w6901 = w48855 ^ w48845;
	assign w6983 = w28752 ^ w48848;
	assign w6937 = w7152 ^ w48856;
	assign w7222 = w6937 ^ w6938;
	assign w7020 = w48856 ^ w34379;
	assign w47489 = w48730 ^ w1456;
	assign w7150 = w48853 ^ w48858;
	assign w7092 = w7201 ^ w7150;
	assign w48726 = w48842 ^ w7092;
	assign w47493 = w48726 ^ w1452;
	assign w7074 = w7191 ^ w7150;
	assign w48731 = w7222 ^ w7206;
	assign w47488 = w48731 ^ w1457;
	assign w7195 = w45447 ^ w48857;
	assign w7064 = w7195 ^ w7151;
	assign w7202 = w48852 ^ w48856;
	assign w7095 = w7097 ^ w7202;
	assign w7205 = w48851 ^ w48855;
	assign w7070 = w7206 ^ w7205;
	assign w7068 = ~w7070;
	assign w48722 = w7220 ^ w7205;
	assign w47497 = w48722 ^ w1448;
	assign w7093 = w7203 ^ w7195;
	assign w48725 = w45459 ^ w7093;
	assign w47494 = w48725 ^ w1451;
	assign w7002 = w7195 ^ w45458;
	assign w7077 = w7201 ^ w28752;
	assign w48733 = w7077 ^ w7078;
	assign w47486 = w48733 ^ w1459;
	assign w25178 = w47488 ^ w47486;
	assign w48735 = w45461 ^ w7074;
	assign w47484 = w48735 ^ w1461;
	assign w7067 = w7203 ^ w7202;
	assign w48740 = w45446 ^ w7067;
	assign w47479 = w48740 ^ w1466;
	assign w48742 = w48853 ^ w7064;
	assign w47477 = w48742 ^ w1468;
	assign w31608 = w47479 ^ w47477;
	assign w44572 = w28699 ^ w28701;
	assign w28657 = w44572 ^ w28654;
	assign w28754 = w28656 ^ w28657;
	assign w28644 = w28648 ^ w44572;
	assign w28647 = w28686 ^ w28644;
	assign w28751 = w28646 ^ w28647;
	assign w28643 = w28667 ^ w28644;
	assign w48854 = w28642 ^ w28643;
	assign w7193 = w48839 ^ w48854;
	assign w7055 = ~w7193;
	assign w7052 = w7205 ^ w7055;
	assign w7124 = w7055 ^ w45792;
	assign w48721 = w7124 ^ w7125;
	assign w47498 = w48721 ^ w1447;
	assign w13494 = w47497 ^ w47498;
	assign w13605 = w47493 ^ w47498;
	assign w7087 = w7193 ^ w7192;
	assign w48729 = w48843 ^ w7087;
	assign w47490 = w48729 ^ w1455;
	assign w25266 = w47490 ^ w47488;
	assign w25152 = w47489 ^ w47490;
	assign w7158 = w48842 ^ w48858;
	assign w7054 = ~w7158;
	assign w6900 = w7158 ^ w48840;
	assign w7237 = w6900 ^ w6901;
	assign w48715 = w7237 ^ w7202;
	assign w47504 = w48715 ^ w1441;
	assign w7143 = w7191 ^ w7158;
	assign w7053 = w7054 ^ w48844;
	assign w48714 = w7052 ^ w7053;
	assign w47505 = w48714 ^ w1440;
	assign w7141 = w7170 ^ w7161;
	assign w45558 = ~w25535;
	assign w7123 = w25536 ^ w45558;
	assign w7179 = w45558 ^ w45646;
	assign w7113 = w7179 ^ w48906;
	assign w7137 = w7179 ^ w7167;
	assign w45559 = ~w25537;
	assign w6953 = w7162 ^ w45559;
	assign w45560 = ~w25538;
	assign w6910 = w7156 ^ w45560;
	assign w45651 = ~w28751;
	assign w7079 = w7203 ^ w45651;
	assign w7198 = w45446 ^ w45651;
	assign w7065 = w7201 ^ w7198;
	assign w48741 = w45447 ^ w7065;
	assign w7021 = w7198 ^ w48841;
	assign w7019 = ~w7021;
	assign w48716 = w7019 ^ w7020;
	assign w47478 = w48741 ^ w1467;
	assign w31614 = w47484 ^ w47478;
	assign w31691 = w31608 ^ w31614;
	assign w31694 = w47479 ^ w31614;
	assign w47503 = w48716 ^ w1442;
	assign w7094 = w7206 ^ w7198;
	assign w48724 = w45458 ^ w7094;
	assign w47495 = w48724 ^ w1450;
	assign w13518 = w47495 ^ w47493;
	assign w48732 = w7079 ^ w7080;
	assign w47487 = w48732 ^ w1458;
	assign w25137 = w25178 ^ w47487;
	assign w7003 = w45651 ^ w34380;
	assign w7001 = w7002 ^ w7003;
	assign w48717 = ~w7001;
	assign w47502 = w48717 ^ w1443;
	assign w19952 = w47504 ^ w47502;
	assign w19911 = w19952 ^ w47503;
	assign w45652 = ~w28753;
	assign w7083 = w7054 ^ w45652;
	assign w7213 = w45460 ^ w45652;
	assign w7089 = w7213 ^ w7191;
	assign w7066 = w7213 ^ w7190;
	assign w48713 = w48854 ^ w7066;
	assign w7088 = w7089 ^ w7090;
	assign w47506 = w48713 ^ w1439;
	assign w20040 = w47506 ^ w47504;
	assign w19926 = w47505 ^ w47506;
	assign w48728 = ~w7088;
	assign w47491 = w48728 ^ w1454;
	assign w25175 = w47491 ^ w47489;
	assign w25177 = w47490 ^ w25175;
	assign w25253 = w47486 ^ w25177;
	assign w25250 = w47487 ^ w25177;
	assign w25192 = w47491 ^ w47490;
	assign w7072 = w45652 ^ w20177;
	assign w48737 = w7071 ^ w7072;
	assign w47482 = w48737 ^ w1463;
	assign w31695 = w47477 ^ w47482;
	assign w45653 = ~w28754;
	assign w6943 = w7150 ^ w45653;
	assign w7219 = w6943 ^ w6944;
	assign w48736 = w7219 ^ w7192;
	assign w47483 = w48736 ^ w1462;
	assign w31690 = w47483 ^ w31694;
	assign w31624 = w47483 ^ w47482;
	assign w31689 = w31624 ^ w31691;
	assign w31697 = w47477 ^ w47483;
	assign w31677 = w31694 & w31690;
	assign w7214 = w45461 ^ w45653;
	assign w7091 = w7214 ^ w7152;
	assign w48727 = w45793 ^ w7091;
	assign w7082 = w7214 ^ w7192;
	assign w6966 = w7214 ^ w7151;
	assign w48719 = w45448 ^ w6966;
	assign w7081 = w7082 ^ w7083;
	assign w48712 = ~w7081;
	assign w47507 = w48712 ^ w1438;
	assign w19949 = w47507 ^ w47505;
	assign w19951 = w47506 ^ w19949;
	assign w20027 = w47502 ^ w19951;
	assign w20024 = w47503 ^ w19951;
	assign w19966 = w47507 ^ w47506;
	assign w47500 = w48719 ^ w1445;
	assign w13524 = w47500 ^ w47494;
	assign w13601 = w13518 ^ w13524;
	assign w13604 = w47495 ^ w13524;
	assign w48711 = w45653 ^ w7143;
	assign w47508 = w48711 ^ w1437;
	assign w19956 = w47508 ^ w47502;
	assign w20026 = w19956 ^ w19951;
	assign w20036 = w47503 ^ w19956;
	assign w20032 = w47507 ^ w20036;
	assign w20035 = w47508 ^ w19911;
	assign w20021 = w47508 & w20035;
	assign w20019 = w20036 & w20032;
	assign w47492 = w48727 ^ w1453;
	assign w25182 = w47492 ^ w47486;
	assign w25252 = w25182 ^ w25177;
	assign w25262 = w47487 ^ w25182;
	assign w25258 = w47491 ^ w25262;
	assign w25261 = w47492 ^ w25137;
	assign w25247 = w47492 & w25261;
	assign w25245 = w25262 & w25258;
	assign w45909 = ~w6669;
	assign w6567 = w45909 ^ w48659;
	assign w48553 = w6566 ^ w6567;
	assign w6564 = w45909 ^ w48660;
	assign w48554 = w6563 ^ w6564;
	assign w47592 = w48554 ^ w1958;
	assign w13788 = w47592 ^ w47590;
	assign w13874 = w47592 ^ w47589;
	assign w13876 = w47594 ^ w47592;
	assign w13861 = w13786 ^ w13876;
	assign w13748 = w13788 ^ w13786;
	assign w13747 = w13788 ^ w47591;
	assign w13871 = w47596 ^ w13747;
	assign w13857 = w47596 & w13871;
	assign w13852 = w13876 & w13861;
	assign w6571 = w45909 ^ w45477;
	assign w6569 = w6570 ^ w6571;
	assign w47593 = w48553 ^ w1957;
	assign w13762 = w47593 ^ w47594;
	assign w48551 = ~w6569;
	assign w47595 = w48551 ^ w1955;
	assign w13875 = w47589 ^ w47595;
	assign w13785 = w47595 ^ w47593;
	assign w13787 = w47594 ^ w13785;
	assign w13860 = w47591 ^ w13787;
	assign w13863 = w47590 ^ w13787;
	assign w13862 = w13792 ^ w13787;
	assign w13868 = w47595 ^ w13872;
	assign w13866 = w13785 ^ w13874;
	assign w13865 = w47596 ^ w13866;
	assign w13802 = w47595 ^ w47594;
	assign w13870 = w13874 ^ w13802;
	assign w13867 = w13802 ^ w13869;
	assign w13864 = w13785 ^ w13748;
	assign w13853 = w13874 & w13863;
	assign w13789 = w13853 ^ w13787;
	assign w13859 = w13866 & w13870;
	assign w13791 = w13859 ^ w13788;
	assign w13795 = w13791 ^ w13789;
	assign w13800 = w47589 ^ w13795;
	assign w13858 = w13867 & w13865;
	assign w13809 = w13852 ^ w13858;
	assign w13850 = w13809 ^ w13800;
	assign w13856 = w13875 & w13860;
	assign w13790 = w13856 ^ w13786;
	assign w13855 = w13872 & w13868;
	assign w13854 = w13869 & w13862;
	assign w13851 = w13873 & w13864;
	assign w13761 = w13852 ^ w13853;
	assign w43947 = w13851 ^ w13854;
	assign w13764 = w13790 ^ w43947;
	assign w13848 = w13764 ^ w13789;
	assign w13804 = w13852 ^ w43947;
	assign w13760 = w13855 ^ w13804;
	assign w13842 = w47595 ^ w13760;
	assign w43950 = w13851 ^ w13857;
	assign w13763 = w13795 ^ w43950;
	assign w13806 = w47591 ^ w13763;
	assign w13801 = w43950 ^ w13786;
	assign w13847 = w13809 ^ w13801;
	assign w13808 = w13761 ^ w13762;
	assign w13807 = w13808 ^ w13790;
	assign w13849 = w13855 ^ w13807;
	assign w13846 = w13850 & w13849;
	assign w13845 = w13846 ^ w13848;
	assign w13841 = w13846 ^ w13806;
	assign w13844 = w13847 & w13845;
	assign w13843 = w13844 ^ w13806;
	assign w13752 = w13844 ^ w13800;
	assign w13822 = w13843 & w13862;
	assign w13840 = w13841 & w13842;
	assign w13838 = w13846 ^ w13840;
	assign w13839 = w13840 ^ w13848;
	assign w13758 = w13840 ^ w13857;
	assign w13759 = w13840 ^ w13804;
	assign w13816 = w13839 & w13871;
	assign w13825 = w13839 & w47596;
	assign w13837 = w13848 & w13838;
	assign w13835 = w13837 ^ w13845;
	assign w13813 = w13843 & w13869;
	assign w13753 = w13758 ^ w13854;
	assign w13834 = w13843 & w13835;
	assign w13799 = w13834 ^ w13809;
	assign w13833 = w13799 ^ w13801;
	assign w13757 = w13834 ^ w13858;
	assign w13830 = w13799 ^ w13752;
	assign w13823 = w13833 & w13872;
	assign w13815 = w13830 & w13875;
	assign w13814 = w13833 & w13868;
	assign w13784 = w13822 ^ w13814;
	assign w13766 = w13822 ^ w13823;
	assign w13824 = w13830 & w13860;
	assign w13782 = w13824 ^ w13815;
	assign w43949 = w13837 ^ w13855;
	assign w13829 = w43949 ^ w13807;
	assign w13827 = w13829 & w13866;
	assign w13818 = w13829 & w13870;
	assign w13796 = w47595 ^ w43949;
	assign w43951 = w13823 ^ w13824;
	assign w43952 = w13825 ^ w13827;
	assign w13836 = w13796 ^ w13759;
	assign w13817 = w13836 & w13867;
	assign w13826 = w13836 & w13865;
	assign w13749 = w13796 ^ w13757;
	assign w13756 = w13786 ^ w13749;
	assign w13832 = w13753 ^ w13756;
	assign w13810 = w13832 & w13873;
	assign w13819 = w13832 & w13864;
	assign w13797 = w13815 ^ w13819;
	assign w13775 = ~w13797;
	assign w13774 = w13775 ^ w13813;
	assign w13770 = w13774 ^ w43952;
	assign w13755 = w13844 ^ w13856;
	assign w13751 = w13755 ^ w13791;
	assign w13750 = w47591 ^ w13751;
	assign w13828 = w13749 ^ w13750;
	assign w13811 = w13828 & w13876;
	assign w13820 = w13828 & w13861;
	assign w13781 = w13820 ^ w13823;
	assign w13778 = ~w13781;
	assign w13805 = w13820 ^ w43951;
	assign w13771 = w13816 ^ w13805;
	assign w13768 = ~w13771;
	assign w13754 = w47589 ^ w13751;
	assign w13831 = w13753 ^ w13754;
	assign w13821 = w13831 & w13863;
	assign w13777 = w13820 ^ w13821;
	assign w13776 = w13821 ^ w13810;
	assign w13772 = ~w13776;
	assign w13812 = w13831 & w13874;
	assign w13773 = w13812 ^ w13770;
	assign w13877 = w13772 ^ w13773;
	assign w43948 = w13811 ^ w13812;
	assign w13793 = w13817 ^ w43948;
	assign w13769 = w13793 ^ w13770;
	assign w48900 = w13768 ^ w13769;
	assign w6954 = w45648 ^ w48900;
	assign w48809 = w6953 ^ w6954;
	assign w47410 = w48809 ^ w2012;
	assign w7184 = w48895 ^ w48900;
	assign w7105 = w7184 ^ w7174;
	assign w48833 = w48904 ^ w7105;
	assign w47386 = w48833 ^ w2036;
	assign w7117 = w7184 ^ w48908;
	assign w7129 = w7184 ^ w7170;
	assign w7127 = ~w7129;
	assign w13794 = w13818 ^ w13793;
	assign w13798 = w13826 ^ w13794;
	assign w13803 = w13827 ^ w13798;
	assign w48902 = w43951 ^ w13803;
	assign w13878 = w13803 ^ w13777;
	assign w13767 = w13825 ^ w13798;
	assign w48901 = w13766 ^ w13767;
	assign w7164 = w48901 ^ w48905;
	assign w48810 = w7232 ^ w7164;
	assign w7103 = w7164 ^ w7162;
	assign w6899 = w48901 ^ w48900;
	assign w7210 = w48897 ^ w48902;
	assign w7115 = w7210 ^ w7164;
	assign w48835 = w7216 ^ w7210;
	assign w47384 = w48835 ^ w2038;
	assign w31430 = w47386 ^ w47384;
	assign w7126 = w7210 ^ w7179;
	assign w48820 = w45450 ^ w7126;
	assign w47399 = w48820 ^ w2023;
	assign w6949 = w48901 ^ w6950;
	assign w13780 = w13784 ^ w43948;
	assign w13779 = w13775 ^ w13780;
	assign w13783 = w43952 ^ w13780;
	assign w13880 = w13782 ^ w13783;
	assign w13879 = w13778 ^ w13779;
	assign w13765 = w13821 ^ w13805;
	assign w48903 = w13794 ^ w13765;
	assign w7159 = w48903 ^ w48907;
	assign w7116 = w7159 ^ w48910;
	assign w48827 = w7115 ^ w7116;
	assign w47392 = w48827 ^ w2030;
	assign w6896 = w7159 ^ w45648;
	assign w6898 = w7159 ^ w48904;
	assign w7238 = w6898 ^ w6899;
	assign w48826 = w7238 ^ w7170;
	assign w47393 = w48826 ^ w2029;
	assign w7145 = w48899 ^ w48903;
	assign w7098 = w7167 ^ w7145;
	assign w48838 = w48907 ^ w7098;
	assign w47381 = w48838 ^ w2041;
	assign w31428 = w47384 ^ w47381;
	assign w31427 = w47381 ^ w47386;
	assign w7110 = w7145 ^ w48911;
	assign w7136 = w48903 ^ w25536;
	assign w7134 = w7194 ^ w7145;
	assign w48815 = w45560 ^ w7134;
	assign w47404 = w48815 ^ w2018;
	assign w47409 = w48810 ^ w2013;
	assign w19390 = w47409 ^ w47410;
	assign w7142 = w7156 ^ w48902;
	assign w48811 = w7141 ^ w7142;
	assign w47408 = w48811 ^ w2014;
	assign w19504 = w47410 ^ w47408;
	assign w45270 = ~w13880;
	assign w6897 = w45453 ^ w45270;
	assign w7239 = w6896 ^ w6897;
	assign w48807 = w45270 ^ w6955;
	assign w47412 = w48807 ^ w2010;
	assign w7207 = w45560 ^ w45270;
	assign w7119 = w7207 ^ w7159;
	assign w48823 = w45649 ^ w7119;
	assign w7132 = w7207 ^ w7174;
	assign w7109 = w7207 ^ w7144;
	assign w48831 = w45453 ^ w7109;
	assign w47388 = w48831 ^ w2034;
	assign w47396 = w48823 ^ w2026;
	assign w45275 = ~w13877;
	assign w7122 = w7167 ^ w45275;
	assign w7121 = w7122 ^ w7123;
	assign w48821 = ~w7121;
	assign w7114 = w45275 ^ w48902;
	assign w48828 = w7113 ^ w7114;
	assign w47391 = w48828 ^ w2031;
	assign w47398 = w48821 ^ w2024;
	assign w13256 = w47404 ^ w47398;
	assign w13336 = w47399 ^ w13256;
	assign w7169 = w45275 ^ w45450;
	assign w7101 = w7169 ^ w7161;
	assign w48836 = w45558 ^ w7101;
	assign w47383 = w48836 ^ w2039;
	assign w31340 = w47383 ^ w47381;
	assign w31415 = w31340 ^ w31430;
	assign w31406 = w31430 & w31415;
	assign w7140 = ~w7169;
	assign w7138 = w7140 ^ w45646;
	assign w48812 = w7138 ^ w7139;
	assign w47407 = w48812 ^ w2015;
	assign w45276 = ~w13878;
	assign w7111 = w45451 ^ w45276;
	assign w48830 = w7110 ^ w7111;
	assign w47389 = w48830 ^ w2033;
	assign w28258 = w47391 ^ w47389;
	assign w28346 = w47392 ^ w47389;
	assign w48813 = w45276 ^ w7137;
	assign w47406 = w48813 ^ w2016;
	assign w19416 = w47408 ^ w47406;
	assign w19420 = w47412 ^ w47406;
	assign w19500 = w47407 ^ w19420;
	assign w19375 = w19416 ^ w47407;
	assign w19499 = w47412 ^ w19375;
	assign w19485 = w47412 & w19499;
	assign w7209 = w48898 ^ w45276;
	assign w7099 = w7209 ^ w45646;
	assign w7120 = w7209 ^ w7144;
	assign w48837 = w7099 ^ w7100;
	assign w47382 = w48837 ^ w2040;
	assign w31342 = w47384 ^ w47382;
	assign w31346 = w47388 ^ w47382;
	assign w31423 = w31340 ^ w31346;
	assign w31426 = w47383 ^ w31346;
	assign w31302 = w31342 ^ w31340;
	assign w31301 = w31342 ^ w47383;
	assign w31425 = w47388 ^ w31301;
	assign w31411 = w47388 & w31425;
	assign w7112 = w7209 ^ w7169;
	assign w48822 = w48899 ^ w7120;
	assign w48829 = w45647 ^ w7112;
	assign w47390 = w48829 ^ w2032;
	assign w28260 = w47392 ^ w47390;
	assign w28264 = w47396 ^ w47390;
	assign w28341 = w28258 ^ w28264;
	assign w28344 = w47391 ^ w28264;
	assign w28220 = w28260 ^ w28258;
	assign w28219 = w28260 ^ w47391;
	assign w28343 = w47396 ^ w28219;
	assign w28329 = w47396 & w28343;
	assign w47397 = w48822 ^ w2025;
	assign w13250 = w47399 ^ w47397;
	assign w13333 = w13250 ^ w13256;
	assign w45277 = ~w13879;
	assign w6911 = w45649 ^ w45277;
	assign w7233 = w6910 ^ w6911;
	assign w48808 = w7233 ^ w7174;
	assign w47411 = w48808 ^ w2011;
	assign w19413 = w47411 ^ w47409;
	assign w19415 = w47410 ^ w19413;
	assign w19491 = w47406 ^ w19415;
	assign w19488 = w47407 ^ w19415;
	assign w19490 = w19420 ^ w19415;
	assign w19496 = w47411 ^ w19500;
	assign w19430 = w47411 ^ w47410;
	assign w19483 = w19500 & w19496;
	assign w7118 = w45452 ^ w45277;
	assign w48825 = w7117 ^ w7118;
	assign w47394 = w48825 ^ w2028;
	assign w28348 = w47394 ^ w47392;
	assign w28333 = w28258 ^ w28348;
	assign w28234 = w47393 ^ w47394;
	assign w28345 = w47389 ^ w47394;
	assign w28324 = w28348 & w28333;
	assign w7199 = w45559 ^ w45277;
	assign w7108 = ~w7199;
	assign w7106 = w7108 ^ w7194;
	assign w48824 = w7239 ^ w7199;
	assign w47395 = w48824 ^ w2027;
	assign w28257 = w47395 ^ w47393;
	assign w28259 = w47394 ^ w28257;
	assign w28335 = w47390 ^ w28259;
	assign w28332 = w47391 ^ w28259;
	assign w28334 = w28264 ^ w28259;
	assign w28340 = w47395 ^ w28344;
	assign w28338 = w28257 ^ w28346;
	assign w28337 = w47396 ^ w28338;
	assign w28274 = w47395 ^ w47394;
	assign w28339 = w28274 ^ w28341;
	assign w28342 = w28346 ^ w28274;
	assign w28336 = w28257 ^ w28220;
	assign w28347 = w47389 ^ w47395;
	assign w28331 = w28338 & w28342;
	assign w28263 = w28331 ^ w28260;
	assign w28330 = w28339 & w28337;
	assign w28281 = w28324 ^ w28330;
	assign w28328 = w28347 & w28332;
	assign w28262 = w28328 ^ w28258;
	assign w28327 = w28344 & w28340;
	assign w28326 = w28341 & w28334;
	assign w28325 = w28346 & w28335;
	assign w28261 = w28325 ^ w28259;
	assign w28267 = w28263 ^ w28261;
	assign w28272 = w47389 ^ w28267;
	assign w28322 = w28281 ^ w28272;
	assign w28233 = w28324 ^ w28325;
	assign w28280 = w28233 ^ w28234;
	assign w28279 = w28280 ^ w28262;
	assign w28321 = w28327 ^ w28279;
	assign w28323 = w28345 & w28336;
	assign w28318 = w28322 & w28321;
	assign w7130 = w7199 ^ w7162;
	assign w48817 = w48895 ^ w7130;
	assign w47402 = w48817 ^ w2020;
	assign w13337 = w47397 ^ w47402;
	assign w44551 = w28323 ^ w28326;
	assign w28236 = w28262 ^ w44551;
	assign w28320 = w28236 ^ w28261;
	assign w28317 = w28318 ^ w28320;
	assign w28276 = w28324 ^ w44551;
	assign w28232 = w28327 ^ w28276;
	assign w28314 = w47395 ^ w28232;
	assign w44554 = w28323 ^ w28329;
	assign w28235 = w28267 ^ w44554;
	assign w28278 = w47391 ^ w28235;
	assign w28313 = w28318 ^ w28278;
	assign w28312 = w28313 & w28314;
	assign w28310 = w28318 ^ w28312;
	assign w28231 = w28312 ^ w28276;
	assign w28230 = w28312 ^ w28329;
	assign w28225 = w28230 ^ w28326;
	assign w28309 = w28320 & w28310;
	assign w28307 = w28309 ^ w28317;
	assign w44553 = w28309 ^ w28327;
	assign w28301 = w44553 ^ w28279;
	assign w28290 = w28301 & w28342;
	assign w28299 = w28301 & w28338;
	assign w28268 = w47395 ^ w44553;
	assign w28308 = w28268 ^ w28231;
	assign w28298 = w28308 & w28337;
	assign w28289 = w28308 & w28339;
	assign w28311 = w28312 ^ w28320;
	assign w28297 = w28311 & w47396;
	assign w28288 = w28311 & w28343;
	assign w28273 = w44554 ^ w28258;
	assign w28319 = w28281 ^ w28273;
	assign w28316 = w28319 & w28317;
	assign w28315 = w28316 ^ w28278;
	assign w28227 = w28316 ^ w28328;
	assign w28223 = w28227 ^ w28263;
	assign w28226 = w47389 ^ w28223;
	assign w28303 = w28225 ^ w28226;
	assign w28224 = w28316 ^ w28272;
	assign w28222 = w47391 ^ w28223;
	assign w28306 = w28315 & w28307;
	assign w28271 = w28306 ^ w28281;
	assign w28305 = w28271 ^ w28273;
	assign w28229 = w28306 ^ w28330;
	assign w28221 = w28268 ^ w28229;
	assign w28228 = w28258 ^ w28221;
	assign w28304 = w28225 ^ w28228;
	assign w28302 = w28271 ^ w28224;
	assign w28300 = w28221 ^ w28222;
	assign w28296 = w28302 & w28332;
	assign w28295 = w28305 & w28344;
	assign w28294 = w28315 & w28334;
	assign w28238 = w28294 ^ w28295;
	assign w28293 = w28303 & w28335;
	assign w28292 = w28300 & w28333;
	assign w28253 = w28292 ^ w28295;
	assign w28250 = ~w28253;
	assign w28249 = w28292 ^ w28293;
	assign w28291 = w28304 & w28336;
	assign w28287 = w28302 & w28347;
	assign w28269 = w28287 ^ w28291;
	assign w28254 = w28296 ^ w28287;
	assign w28247 = ~w28269;
	assign w28286 = w28305 & w28340;
	assign w28256 = w28294 ^ w28286;
	assign w28285 = w28315 & w28341;
	assign w28246 = w28247 ^ w28285;
	assign w28284 = w28303 & w28346;
	assign w28283 = w28300 & w28348;
	assign w28282 = w28304 & w28345;
	assign w28248 = w28293 ^ w28282;
	assign w28244 = ~w28248;
	assign w44552 = w28283 ^ w28284;
	assign w28265 = w28289 ^ w44552;
	assign w28266 = w28290 ^ w28265;
	assign w28270 = w28298 ^ w28266;
	assign w28239 = w28297 ^ w28270;
	assign w49052 = w28238 ^ w28239;
	assign w7282 = w49052 ^ w49045;
	assign w28275 = w28299 ^ w28270;
	assign w28350 = w28275 ^ w28249;
	assign w28252 = w28256 ^ w44552;
	assign w28251 = w28247 ^ w28252;
	assign w28351 = w28250 ^ w28251;
	assign w49050 = ~w28351;
	assign w7284 = w28351 ^ w45439;
	assign w7536 = w45267 ^ w49050;
	assign w44555 = w28295 ^ w28296;
	assign w49053 = w44555 ^ w28275;
	assign w7424 = w49053 ^ w49046;
	assign w28277 = w28292 ^ w44555;
	assign w28243 = w28288 ^ w28277;
	assign w28240 = ~w28243;
	assign w28237 = w28293 ^ w28277;
	assign w49054 = w28266 ^ w28237;
	assign w7496 = w49049 ^ w49054;
	assign w7430 = ~w7496;
	assign w7434 = w7430 ^ w45267;
	assign w44556 = w28297 ^ w28299;
	assign w28255 = w44556 ^ w28252;
	assign w28352 = w28254 ^ w28255;
	assign w28242 = w28246 ^ w44556;
	assign w28245 = w28284 ^ w28242;
	assign w28349 = w28244 ^ w28245;
	assign w28241 = w28265 ^ w28242;
	assign w49051 = w28240 ^ w28241;
	assign w7534 = w49044 ^ w49051;
	assign w7291 = ~w49051;
	assign w7417 = ~w7534;
	assign w7415 = w7417 ^ w49040;
	assign w7428 = w7559 ^ w7417;
	assign w7290 = w49052 ^ w7291;
	assign w7469 = w45438 ^ w7291;
	assign w45638 = ~w28349;
	assign w7422 = w45638 ^ w13475;
	assign w45639 = ~w28350;
	assign w7420 = w45639 ^ w13476;
	assign w45640 = ~w28352;
	assign w7288 = w45438 ^ w45640;
	assign w7535 = w45268 ^ w45640;
	assign w45910 = ~w7144;
	assign w7107 = w45910 ^ w45452;
	assign w48832 = w7106 ^ w7107;
	assign w47387 = w48832 ^ w2035;
	assign w31422 = w47387 ^ w31426;
	assign w31356 = w47387 ^ w47386;
	assign w31421 = w31356 ^ w31423;
	assign w31424 = w31428 ^ w31356;
	assign w31429 = w47381 ^ w47387;
	assign w31409 = w31426 & w31422;
	assign w7104 = w45910 ^ w48896;
	assign w7102 = w7103 ^ w7104;
	assign w48834 = ~w7102;
	assign w47385 = w48834 ^ w2037;
	assign w31339 = w47387 ^ w47385;
	assign w31341 = w47386 ^ w31339;
	assign w31417 = w47382 ^ w31341;
	assign w31414 = w47383 ^ w31341;
	assign w31416 = w31346 ^ w31341;
	assign w31420 = w31339 ^ w31428;
	assign w31419 = w47388 ^ w31420;
	assign w31316 = w47385 ^ w47386;
	assign w31418 = w31339 ^ w31302;
	assign w31413 = w31420 & w31424;
	assign w31345 = w31413 ^ w31342;
	assign w31412 = w31421 & w31419;
	assign w31363 = w31406 ^ w31412;
	assign w31410 = w31429 & w31414;
	assign w31344 = w31410 ^ w31340;
	assign w31408 = w31423 & w31416;
	assign w31407 = w31428 & w31417;
	assign w31343 = w31407 ^ w31341;
	assign w31349 = w31345 ^ w31343;
	assign w31354 = w47381 ^ w31349;
	assign w31404 = w31363 ^ w31354;
	assign w31315 = w31406 ^ w31407;
	assign w31362 = w31315 ^ w31316;
	assign w31361 = w31362 ^ w31344;
	assign w31403 = w31409 ^ w31361;
	assign w31405 = w31427 & w31418;
	assign w31400 = w31404 & w31403;
	assign w7135 = w45910 ^ w45647;
	assign w48814 = w7135 ^ w7136;
	assign w47405 = w48814 ^ w2017;
	assign w19414 = w47407 ^ w47405;
	assign w19489 = w19414 ^ w19504;
	assign w19502 = w47408 ^ w47405;
	assign w19498 = w19502 ^ w19430;
	assign w19497 = w19414 ^ w19420;
	assign w19495 = w19430 ^ w19497;
	assign w19494 = w19413 ^ w19502;
	assign w19493 = w47412 ^ w19494;
	assign w19376 = w19416 ^ w19414;
	assign w19492 = w19413 ^ w19376;
	assign w19503 = w47405 ^ w47411;
	assign w19501 = w47405 ^ w47410;
	assign w19487 = w19494 & w19498;
	assign w19419 = w19487 ^ w19416;
	assign w19486 = w19495 & w19493;
	assign w19484 = w19503 & w19488;
	assign w19418 = w19484 ^ w19414;
	assign w19482 = w19497 & w19490;
	assign w19481 = w19502 & w19491;
	assign w19417 = w19481 ^ w19415;
	assign w19423 = w19419 ^ w19417;
	assign w19428 = w47405 ^ w19423;
	assign w19480 = w19504 & w19489;
	assign w19437 = w19480 ^ w19486;
	assign w19478 = w19437 ^ w19428;
	assign w19389 = w19480 ^ w19481;
	assign w19436 = w19389 ^ w19390;
	assign w19435 = w19436 ^ w19418;
	assign w19477 = w19483 ^ w19435;
	assign w19479 = w19501 & w19492;
	assign w19474 = w19478 & w19477;
	assign w44182 = w19479 ^ w19482;
	assign w19392 = w19418 ^ w44182;
	assign w19476 = w19392 ^ w19417;
	assign w19473 = w19474 ^ w19476;
	assign w19432 = w19480 ^ w44182;
	assign w19388 = w19483 ^ w19432;
	assign w19470 = w47411 ^ w19388;
	assign w44185 = w19479 ^ w19485;
	assign w19391 = w19423 ^ w44185;
	assign w19434 = w47407 ^ w19391;
	assign w19469 = w19474 ^ w19434;
	assign w19468 = w19469 & w19470;
	assign w19467 = w19468 ^ w19476;
	assign w19466 = w19474 ^ w19468;
	assign w19387 = w19468 ^ w19432;
	assign w19386 = w19468 ^ w19485;
	assign w19381 = w19386 ^ w19482;
	assign w19465 = w19476 & w19466;
	assign w19463 = w19465 ^ w19473;
	assign w19453 = w19467 & w47412;
	assign w19444 = w19467 & w19499;
	assign w44184 = w19465 ^ w19483;
	assign w19457 = w44184 ^ w19435;
	assign w19455 = w19457 & w19494;
	assign w19446 = w19457 & w19498;
	assign w19424 = w47411 ^ w44184;
	assign w19464 = w19424 ^ w19387;
	assign w19454 = w19464 & w19493;
	assign w19445 = w19464 & w19495;
	assign w19429 = w44185 ^ w19414;
	assign w19475 = w19437 ^ w19429;
	assign w19472 = w19475 & w19473;
	assign w19471 = w19472 ^ w19434;
	assign w19383 = w19472 ^ w19484;
	assign w19379 = w19383 ^ w19419;
	assign w19382 = w47405 ^ w19379;
	assign w19459 = w19381 ^ w19382;
	assign w19380 = w19472 ^ w19428;
	assign w19378 = w47407 ^ w19379;
	assign w19462 = w19471 & w19463;
	assign w19427 = w19462 ^ w19437;
	assign w19461 = w19427 ^ w19429;
	assign w19385 = w19462 ^ w19486;
	assign w19377 = w19424 ^ w19385;
	assign w19384 = w19414 ^ w19377;
	assign w19460 = w19381 ^ w19384;
	assign w19458 = w19427 ^ w19380;
	assign w19456 = w19377 ^ w19378;
	assign w19452 = w19458 & w19488;
	assign w19451 = w19461 & w19500;
	assign w19450 = w19471 & w19490;
	assign w19394 = w19450 ^ w19451;
	assign w19449 = w19459 & w19491;
	assign w19448 = w19456 & w19489;
	assign w19409 = w19448 ^ w19451;
	assign w19406 = ~w19409;
	assign w19405 = w19448 ^ w19449;
	assign w19447 = w19460 & w19492;
	assign w19443 = w19458 & w19503;
	assign w19425 = w19443 ^ w19447;
	assign w19410 = w19452 ^ w19443;
	assign w19403 = ~w19425;
	assign w19442 = w19461 & w19496;
	assign w19412 = w19450 ^ w19442;
	assign w19441 = w19471 & w19497;
	assign w19402 = w19403 ^ w19441;
	assign w19440 = w19459 & w19502;
	assign w19439 = w19456 & w19504;
	assign w19438 = w19460 & w19501;
	assign w19404 = w19449 ^ w19438;
	assign w19400 = ~w19404;
	assign w44183 = w19439 ^ w19440;
	assign w19421 = w19445 ^ w44183;
	assign w19422 = w19446 ^ w19421;
	assign w19426 = w19454 ^ w19422;
	assign w19431 = w19455 ^ w19426;
	assign w19506 = w19431 ^ w19405;
	assign w19395 = w19453 ^ w19426;
	assign w49078 = w19394 ^ w19395;
	assign w19408 = w19412 ^ w44183;
	assign w19407 = w19403 ^ w19408;
	assign w19507 = w19406 ^ w19407;
	assign w44186 = w19451 ^ w19452;
	assign w49079 = w44186 ^ w19431;
	assign w19433 = w19448 ^ w44186;
	assign w19399 = w19444 ^ w19433;
	assign w19396 = ~w19399;
	assign w19393 = w19449 ^ w19433;
	assign w49080 = w19422 ^ w19393;
	assign w44187 = w19453 ^ w19455;
	assign w19411 = w44187 ^ w19408;
	assign w19508 = w19410 ^ w19411;
	assign w19398 = w19402 ^ w44187;
	assign w19401 = w19440 ^ w19398;
	assign w19505 = w19400 ^ w19401;
	assign w19397 = w19421 ^ w19398;
	assign w49077 = w19396 ^ w19397;
	assign w44683 = w31405 ^ w31411;
	assign w31355 = w44683 ^ w31340;
	assign w31401 = w31363 ^ w31355;
	assign w31317 = w31349 ^ w44683;
	assign w31360 = w47383 ^ w31317;
	assign w31395 = w31400 ^ w31360;
	assign w44684 = w31405 ^ w31408;
	assign w31358 = w31406 ^ w44684;
	assign w31314 = w31409 ^ w31358;
	assign w31396 = w47387 ^ w31314;
	assign w31394 = w31395 & w31396;
	assign w31313 = w31394 ^ w31358;
	assign w31312 = w31394 ^ w31411;
	assign w31307 = w31312 ^ w31408;
	assign w31392 = w31400 ^ w31394;
	assign w31318 = w31344 ^ w44684;
	assign w31402 = w31318 ^ w31343;
	assign w31393 = w31394 ^ w31402;
	assign w31399 = w31400 ^ w31402;
	assign w31398 = w31401 & w31399;
	assign w31397 = w31398 ^ w31360;
	assign w31309 = w31398 ^ w31410;
	assign w31305 = w31309 ^ w31345;
	assign w31308 = w47381 ^ w31305;
	assign w31385 = w31307 ^ w31308;
	assign w31306 = w31398 ^ w31354;
	assign w31304 = w47383 ^ w31305;
	assign w31391 = w31402 & w31392;
	assign w31389 = w31391 ^ w31399;
	assign w31388 = w31397 & w31389;
	assign w31353 = w31388 ^ w31363;
	assign w31387 = w31353 ^ w31355;
	assign w31311 = w31388 ^ w31412;
	assign w31384 = w31353 ^ w31306;
	assign w31379 = w31393 & w47388;
	assign w31378 = w31384 & w31414;
	assign w31377 = w31387 & w31426;
	assign w31376 = w31397 & w31416;
	assign w31320 = w31376 ^ w31377;
	assign w31375 = w31385 & w31417;
	assign w31370 = w31393 & w31425;
	assign w31369 = w31384 & w31429;
	assign w31336 = w31378 ^ w31369;
	assign w31368 = w31387 & w31422;
	assign w31338 = w31376 ^ w31368;
	assign w31367 = w31397 & w31423;
	assign w31366 = w31385 & w31428;
	assign w44685 = w31377 ^ w31378;
	assign w44687 = w31391 ^ w31409;
	assign w31350 = w47387 ^ w44687;
	assign w31390 = w31350 ^ w31313;
	assign w31371 = w31390 & w31421;
	assign w31380 = w31390 & w31419;
	assign w31303 = w31350 ^ w31311;
	assign w31310 = w31340 ^ w31303;
	assign w31386 = w31307 ^ w31310;
	assign w31373 = w31386 & w31418;
	assign w31351 = w31369 ^ w31373;
	assign w31329 = ~w31351;
	assign w31328 = w31329 ^ w31367;
	assign w31382 = w31303 ^ w31304;
	assign w31365 = w31382 & w31430;
	assign w31364 = w31386 & w31427;
	assign w31330 = w31375 ^ w31364;
	assign w31326 = ~w31330;
	assign w43586 = w31365 ^ w31366;
	assign w31347 = w31371 ^ w43586;
	assign w31334 = w31338 ^ w43586;
	assign w31333 = w31329 ^ w31334;
	assign w31374 = w31382 & w31415;
	assign w31331 = w31374 ^ w31375;
	assign w31359 = w31374 ^ w44685;
	assign w31325 = w31370 ^ w31359;
	assign w31322 = ~w31325;
	assign w31319 = w31375 ^ w31359;
	assign w31335 = w31374 ^ w31377;
	assign w31332 = ~w31335;
	assign w31433 = w31332 ^ w31333;
	assign w31383 = w44687 ^ w31361;
	assign w31381 = w31383 & w31420;
	assign w31372 = w31383 & w31424;
	assign w31348 = w31372 ^ w31347;
	assign w31352 = w31380 ^ w31348;
	assign w31357 = w31381 ^ w31352;
	assign w49111 = w44685 ^ w31357;
	assign w31432 = w31357 ^ w31331;
	assign w31321 = w31379 ^ w31352;
	assign w49110 = w31320 ^ w31321;
	assign w49112 = w31348 ^ w31319;
	assign w7488 = w49108 ^ w49112;
	assign w7505 = w49107 ^ w49111;
	assign w7295 = w7488 ^ w49110;
	assign w7560 = w7295 ^ w7296;
	assign w44686 = w31379 ^ w31381;
	assign w31337 = w44686 ^ w31334;
	assign w31434 = w31336 ^ w31337;
	assign w31324 = w31328 ^ w44686;
	assign w31327 = w31366 ^ w31324;
	assign w31431 = w31326 ^ w31327;
	assign w31323 = w31347 ^ w31324;
	assign w49109 = w31322 ^ w31323;
	assign w7506 = w49105 ^ w49109;
	assign w7257 = w49110 ^ w49109;
	assign w45426 = ~w19507;
	assign w45427 = ~w19508;
	assign w45432 = ~w19505;
	assign w45433 = ~w19506;
	assign w45722 = ~w31432;
	assign w7511 = w45437 ^ w45722;
	assign w45723 = ~w31433;
	assign w7518 = w45430 ^ w45723;
	assign w45724 = ~w31434;
	assign w7538 = w45431 ^ w45724;
	assign w45729 = ~w31431;
	assign w45911 = ~w7150;
	assign w6945 = w45911 ^ w48854;
	assign w6982 = w45911 ^ w45459;
	assign w7218 = w6945 ^ w6946;
	assign w48718 = w6982 ^ w6983;
	assign w7069 = w45911 ^ w48852;
	assign w47501 = w48718 ^ w1444;
	assign w19950 = w47503 ^ w47501;
	assign w20025 = w19950 ^ w20040;
	assign w20038 = w47504 ^ w47501;
	assign w20034 = w20038 ^ w19966;
	assign w20033 = w19950 ^ w19956;
	assign w20031 = w19966 ^ w20033;
	assign w20030 = w19949 ^ w20038;
	assign w20029 = w47508 ^ w20030;
	assign w19912 = w19952 ^ w19950;
	assign w20028 = w19949 ^ w19912;
	assign w20039 = w47501 ^ w47507;
	assign w20037 = w47501 ^ w47506;
	assign w20023 = w20030 & w20034;
	assign w19955 = w20023 ^ w19952;
	assign w20022 = w20031 & w20029;
	assign w20020 = w20039 & w20024;
	assign w19954 = w20020 ^ w19950;
	assign w20018 = w20033 & w20026;
	assign w20017 = w20038 & w20027;
	assign w19953 = w20017 ^ w19951;
	assign w19959 = w19955 ^ w19953;
	assign w19964 = w47501 ^ w19959;
	assign w20016 = w20040 & w20025;
	assign w19973 = w20016 ^ w20022;
	assign w20014 = w19973 ^ w19964;
	assign w19925 = w20016 ^ w20017;
	assign w19972 = w19925 ^ w19926;
	assign w19971 = w19972 ^ w19954;
	assign w20013 = w20019 ^ w19971;
	assign w20015 = w20037 & w20028;
	assign w20010 = w20014 & w20013;
	assign w48738 = w7218 ^ w7215;
	assign w47481 = w48738 ^ w1464;
	assign w31607 = w47483 ^ w47481;
	assign w31609 = w47482 ^ w31607;
	assign w31685 = w47478 ^ w31609;
	assign w31682 = w47479 ^ w31609;
	assign w31684 = w31614 ^ w31609;
	assign w31584 = w47481 ^ w47482;
	assign w31678 = w31697 & w31682;
	assign w31612 = w31678 ^ w31608;
	assign w31676 = w31691 & w31684;
	assign w48739 = w7068 ^ w7069;
	assign w47480 = w48739 ^ w1465;
	assign w31610 = w47480 ^ w47478;
	assign w31696 = w47480 ^ w47477;
	assign w31692 = w31696 ^ w31624;
	assign w31688 = w31607 ^ w31696;
	assign w31687 = w47484 ^ w31688;
	assign w31698 = w47482 ^ w47480;
	assign w31683 = w31608 ^ w31698;
	assign w31570 = w31610 ^ w31608;
	assign w31686 = w31607 ^ w31570;
	assign w31569 = w31610 ^ w47479;
	assign w31693 = w47484 ^ w31569;
	assign w31681 = w31688 & w31692;
	assign w31613 = w31681 ^ w31610;
	assign w31680 = w31689 & w31687;
	assign w31679 = w47484 & w31693;
	assign w31675 = w31696 & w31685;
	assign w31611 = w31675 ^ w31609;
	assign w31617 = w31613 ^ w31611;
	assign w31622 = w47477 ^ w31617;
	assign w31674 = w31698 & w31683;
	assign w31631 = w31674 ^ w31680;
	assign w31672 = w31631 ^ w31622;
	assign w31583 = w31674 ^ w31675;
	assign w31630 = w31583 ^ w31584;
	assign w31629 = w31630 ^ w31612;
	assign w31671 = w31677 ^ w31629;
	assign w31673 = w31695 & w31686;
	assign w31668 = w31672 & w31671;
	assign w44205 = w20015 ^ w20021;
	assign w19927 = w19959 ^ w44205;
	assign w19970 = w47503 ^ w19927;
	assign w20005 = w20010 ^ w19970;
	assign w19965 = w44205 ^ w19950;
	assign w20011 = w19973 ^ w19965;
	assign w44206 = w20015 ^ w20018;
	assign w19968 = w20016 ^ w44206;
	assign w19924 = w20019 ^ w19968;
	assign w20006 = w47507 ^ w19924;
	assign w20004 = w20005 & w20006;
	assign w19923 = w20004 ^ w19968;
	assign w19922 = w20004 ^ w20021;
	assign w20002 = w20010 ^ w20004;
	assign w19917 = w19922 ^ w20018;
	assign w19928 = w19954 ^ w44206;
	assign w20012 = w19928 ^ w19953;
	assign w20003 = w20004 ^ w20012;
	assign w20009 = w20010 ^ w20012;
	assign w20008 = w20011 & w20009;
	assign w20007 = w20008 ^ w19970;
	assign w19919 = w20008 ^ w20020;
	assign w19915 = w19919 ^ w19955;
	assign w19918 = w47501 ^ w19915;
	assign w19995 = w19917 ^ w19918;
	assign w19916 = w20008 ^ w19964;
	assign w19914 = w47503 ^ w19915;
	assign w20001 = w20012 & w20002;
	assign w19999 = w20001 ^ w20009;
	assign w19998 = w20007 & w19999;
	assign w19963 = w19998 ^ w19973;
	assign w19997 = w19963 ^ w19965;
	assign w19921 = w19998 ^ w20022;
	assign w19994 = w19963 ^ w19916;
	assign w19989 = w20003 & w47508;
	assign w19988 = w19994 & w20024;
	assign w19987 = w19997 & w20036;
	assign w19986 = w20007 & w20026;
	assign w19930 = w19986 ^ w19987;
	assign w19985 = w19995 & w20027;
	assign w19980 = w20003 & w20035;
	assign w19979 = w19994 & w20039;
	assign w19946 = w19988 ^ w19979;
	assign w19978 = w19997 & w20032;
	assign w19948 = w19986 ^ w19978;
	assign w19977 = w20007 & w20033;
	assign w19976 = w19995 & w20038;
	assign w44207 = w19987 ^ w19988;
	assign w44209 = w20001 ^ w20019;
	assign w19993 = w44209 ^ w19971;
	assign w19991 = w19993 & w20030;
	assign w44208 = w19989 ^ w19991;
	assign w19982 = w19993 & w20034;
	assign w19960 = w47507 ^ w44209;
	assign w20000 = w19960 ^ w19923;
	assign w19913 = w19960 ^ w19921;
	assign w19920 = w19950 ^ w19913;
	assign w19996 = w19917 ^ w19920;
	assign w19992 = w19913 ^ w19914;
	assign w19990 = w20000 & w20029;
	assign w19984 = w19992 & w20025;
	assign w19969 = w19984 ^ w44207;
	assign w19945 = w19984 ^ w19987;
	assign w19942 = ~w19945;
	assign w19941 = w19984 ^ w19985;
	assign w19935 = w19980 ^ w19969;
	assign w19932 = ~w19935;
	assign w19929 = w19985 ^ w19969;
	assign w19983 = w19996 & w20028;
	assign w19961 = w19979 ^ w19983;
	assign w19939 = ~w19961;
	assign w19938 = w19939 ^ w19977;
	assign w19934 = w19938 ^ w44208;
	assign w19937 = w19976 ^ w19934;
	assign w19981 = w20000 & w20031;
	assign w19975 = w19992 & w20040;
	assign w19974 = w19996 & w20037;
	assign w19940 = w19985 ^ w19974;
	assign w19936 = ~w19940;
	assign w20041 = w19936 ^ w19937;
	assign w43554 = w19975 ^ w19976;
	assign w19957 = w19981 ^ w43554;
	assign w19958 = w19982 ^ w19957;
	assign w19962 = w19990 ^ w19958;
	assign w19967 = w19991 ^ w19962;
	assign w49098 = w44207 ^ w19967;
	assign w20042 = w19967 ^ w19941;
	assign w19933 = w19957 ^ w19934;
	assign w49096 = w19932 ^ w19933;
	assign w19931 = w19989 ^ w19962;
	assign w49097 = w19930 ^ w19931;
	assign w49100 = w19958 ^ w19929;
	assign w49099 = ~w20042;
	assign w7500 = w49100 ^ w49112;
	assign w7256 = w7500 ^ w49096;
	assign w7576 = w7256 ^ w7257;
	assign w7294 = ~w49098;
	assign w7483 = w49111 ^ w7294;
	assign w7299 = w7538 ^ w7500;
	assign w19944 = w19948 ^ w43554;
	assign w19947 = w44208 ^ w19944;
	assign w20044 = w19946 ^ w19947;
	assign w19943 = w19939 ^ w19944;
	assign w20043 = w19942 ^ w19943;
	assign w44694 = w31673 ^ w31676;
	assign w31586 = w31612 ^ w44694;
	assign w31670 = w31586 ^ w31611;
	assign w31667 = w31668 ^ w31670;
	assign w31626 = w31674 ^ w44694;
	assign w31582 = w31677 ^ w31626;
	assign w31664 = w47483 ^ w31582;
	assign w44697 = w31673 ^ w31679;
	assign w31585 = w31617 ^ w44697;
	assign w31628 = w47479 ^ w31585;
	assign w31663 = w31668 ^ w31628;
	assign w31662 = w31663 & w31664;
	assign w31660 = w31668 ^ w31662;
	assign w31581 = w31662 ^ w31626;
	assign w31580 = w31662 ^ w31679;
	assign w31575 = w31580 ^ w31676;
	assign w31659 = w31670 & w31660;
	assign w31657 = w31659 ^ w31667;
	assign w44696 = w31659 ^ w31677;
	assign w31651 = w44696 ^ w31629;
	assign w31640 = w31651 & w31692;
	assign w31649 = w31651 & w31688;
	assign w31618 = w47483 ^ w44696;
	assign w31658 = w31618 ^ w31581;
	assign w31648 = w31658 & w31687;
	assign w31639 = w31658 & w31689;
	assign w31661 = w31662 ^ w31670;
	assign w31647 = w31661 & w47484;
	assign w31638 = w31661 & w31693;
	assign w31623 = w44697 ^ w31608;
	assign w31669 = w31631 ^ w31623;
	assign w31666 = w31669 & w31667;
	assign w31665 = w31666 ^ w31628;
	assign w31577 = w31666 ^ w31678;
	assign w31573 = w31577 ^ w31613;
	assign w31576 = w47477 ^ w31573;
	assign w31653 = w31575 ^ w31576;
	assign w31574 = w31666 ^ w31622;
	assign w31572 = w47479 ^ w31573;
	assign w31656 = w31665 & w31657;
	assign w31621 = w31656 ^ w31631;
	assign w31655 = w31621 ^ w31623;
	assign w31579 = w31656 ^ w31680;
	assign w31571 = w31618 ^ w31579;
	assign w31578 = w31608 ^ w31571;
	assign w31654 = w31575 ^ w31578;
	assign w31652 = w31621 ^ w31574;
	assign w31650 = w31571 ^ w31572;
	assign w31646 = w31652 & w31682;
	assign w31645 = w31655 & w31694;
	assign w31644 = w31665 & w31684;
	assign w31588 = w31644 ^ w31645;
	assign w31643 = w31653 & w31685;
	assign w31642 = w31650 & w31683;
	assign w31603 = w31642 ^ w31645;
	assign w31600 = ~w31603;
	assign w31599 = w31642 ^ w31643;
	assign w31641 = w31654 & w31686;
	assign w31637 = w31652 & w31697;
	assign w31619 = w31637 ^ w31641;
	assign w31604 = w31646 ^ w31637;
	assign w31597 = ~w31619;
	assign w31636 = w31655 & w31690;
	assign w31606 = w31644 ^ w31636;
	assign w31635 = w31665 & w31691;
	assign w31596 = w31597 ^ w31635;
	assign w31634 = w31653 & w31696;
	assign w31633 = w31650 & w31698;
	assign w31632 = w31654 & w31695;
	assign w31598 = w31643 ^ w31632;
	assign w31594 = ~w31598;
	assign w44695 = w31633 ^ w31634;
	assign w31615 = w31639 ^ w44695;
	assign w31616 = w31640 ^ w31615;
	assign w31620 = w31648 ^ w31616;
	assign w31589 = w31647 ^ w31620;
	assign w49056 = w31588 ^ w31589;
	assign w7245 = w49056 ^ w49046;
	assign w7549 = w49052 ^ w49056;
	assign w7414 = w7550 ^ w7549;
	assign w48923 = w7564 ^ w7549;
	assign w7429 = w7430 ^ w49056;
	assign w48931 = w7428 ^ w7429;
	assign w47361 = w48931 ^ w1583;
	assign w7412 = ~w7414;
	assign w31625 = w31649 ^ w31620;
	assign w31700 = w31625 ^ w31599;
	assign w49058 = ~w31700;
	assign w7539 = w45639 ^ w49058;
	assign w7346 = w7539 ^ w45444;
	assign w7327 = w31700 ^ w49049;
	assign w7421 = w7545 ^ w31700;
	assign w48934 = w7421 ^ w7422;
	assign w47358 = w48934 ^ w1586;
	assign w7437 = w7547 ^ w7539;
	assign w48926 = w45445 ^ w7437;
	assign w47366 = w48926 ^ w1578;
	assign w7408 = w7539 ^ w7495;
	assign w31602 = w31606 ^ w44695;
	assign w31601 = w31597 ^ w31602;
	assign w31701 = w31600 ^ w31601;
	assign w44698 = w31645 ^ w31646;
	assign w49057 = w44698 ^ w31625;
	assign w7281 = w7496 ^ w49057;
	assign w7566 = w7281 ^ w7282;
	assign w48932 = w7566 ^ w7550;
	assign w47360 = w48932 ^ w1584;
	assign w19148 = w47360 ^ w47358;
	assign w7546 = w49053 ^ w49057;
	assign w7439 = w7441 ^ w7546;
	assign w7411 = w7547 ^ w7546;
	assign w48941 = w45638 ^ w7411;
	assign w47351 = w48941 ^ w1593;
	assign w7364 = w49057 ^ w13475;
	assign w31627 = w31642 ^ w44698;
	assign w31593 = w31638 ^ w31627;
	assign w31590 = ~w31593;
	assign w31587 = w31643 ^ w31627;
	assign w49059 = w31616 ^ w31587;
	assign w7502 = w49043 ^ w49059;
	assign w7494 = w49054 ^ w49059;
	assign w7487 = w7535 ^ w7502;
	assign w7398 = ~w7502;
	assign w7397 = w7398 ^ w49045;
	assign w7418 = w7535 ^ w7494;
	assign w7436 = w7545 ^ w7494;
	assign w48927 = w49043 ^ w7436;
	assign w47365 = w48927 ^ w1579;
	assign w48936 = w45439 ^ w7418;
	assign w47356 = w48936 ^ w1588;
	assign w7244 = w7502 ^ w49041;
	assign w7581 = w7244 ^ w7245;
	assign w48916 = w7581 ^ w7546;
	assign w47376 = w48916 ^ w1568;
	assign w44699 = w31647 ^ w31649;
	assign w31605 = w44699 ^ w31602;
	assign w31702 = w31604 ^ w31605;
	assign w31592 = w31596 ^ w44699;
	assign w31595 = w31634 ^ w31592;
	assign w31699 = w31594 ^ w31595;
	assign w31591 = w31615 ^ w31592;
	assign w49055 = w31590 ^ w31591;
	assign w7537 = w49040 ^ w49055;
	assign w7399 = ~w7537;
	assign w7468 = w7399 ^ w45267;
	assign w48922 = w7468 ^ w7469;
	assign w47370 = w48922 ^ w1574;
	assign w33839 = w47365 ^ w47370;
	assign w7396 = w7549 ^ w7399;
	assign w48915 = w7396 ^ w7397;
	assign w7431 = w7537 ^ w7536;
	assign w48930 = w49044 ^ w7431;
	assign w47362 = w48930 ^ w1582;
	assign w19236 = w47362 ^ w47360;
	assign w19122 = w47361 ^ w47362;
	assign w47377 = w48915 ^ w1567;
	assign w7514 = w49097 ^ w49110;
	assign w7485 = w7514 ^ w7505;
	assign w48943 = w49054 ^ w7408;
	assign w47349 = w48943 ^ w1595;
	assign w31206 = w47351 ^ w47349;
	assign w47369 = w48923 ^ w1575;
	assign w33728 = w47369 ^ w47370;
	assign w45442 = ~w20043;
	assign w7297 = w7506 ^ w45442;
	assign w45443 = ~w20044;
	assign w7254 = w7500 ^ w45443;
	assign w45449 = ~w20041;
	assign w7467 = w20042 ^ w45449;
	assign w7523 = w45449 ^ w45729;
	assign w7481 = w7523 ^ w7511;
	assign w7457 = w7523 ^ w49107;
	assign w45730 = ~w31699;
	assign w7542 = w45638 ^ w45730;
	assign w7365 = w7542 ^ w49042;
	assign w7409 = w7545 ^ w7542;
	assign w48942 = w45639 ^ w7409;
	assign w47350 = w48942 ^ w1594;
	assign w31212 = w47356 ^ w47350;
	assign w31289 = w31206 ^ w31212;
	assign w31292 = w47351 ^ w31212;
	assign w7363 = ~w7365;
	assign w7423 = w7547 ^ w45730;
	assign w7438 = w7550 ^ w7542;
	assign w48925 = w45444 ^ w7438;
	assign w47367 = w48925 ^ w1577;
	assign w33752 = w47367 ^ w47365;
	assign w48933 = w7423 ^ w7424;
	assign w47359 = w48933 ^ w1585;
	assign w19107 = w19148 ^ w47359;
	assign w48917 = w7363 ^ w7364;
	assign w47375 = w48917 ^ w1569;
	assign w7347 = w45730 ^ w13476;
	assign w7345 = w7346 ^ w7347;
	assign w48918 = ~w7345;
	assign w47374 = w48918 ^ w1570;
	assign w19282 = w47376 ^ w47374;
	assign w19241 = w19282 ^ w47375;
	assign w45731 = ~w31701;
	assign w7416 = w45731 ^ w28351;
	assign w48938 = w7415 ^ w7416;
	assign w47354 = w48938 ^ w1590;
	assign w31293 = w47349 ^ w47354;
	assign w7557 = w45438 ^ w45731;
	assign w7410 = w7557 ^ w7534;
	assign w7433 = w7557 ^ w7535;
	assign w7432 = w7433 ^ w7434;
	assign w48929 = ~w7432;
	assign w47363 = w48929 ^ w1581;
	assign w19145 = w47363 ^ w47361;
	assign w19147 = w47362 ^ w19145;
	assign w19223 = w47358 ^ w19147;
	assign w19220 = w47359 ^ w19147;
	assign w19162 = w47363 ^ w47362;
	assign w7427 = w7398 ^ w45731;
	assign w48914 = w49055 ^ w7410;
	assign w47378 = w48914 ^ w1566;
	assign w19370 = w47378 ^ w47376;
	assign w19256 = w47377 ^ w47378;
	assign w45732 = ~w31702;
	assign w7287 = w7494 ^ w45732;
	assign w7563 = w7287 ^ w7288;
	assign w48937 = w7563 ^ w7536;
	assign w7558 = w45439 ^ w45732;
	assign w48912 = w45732 ^ w7487;
	assign w7310 = w7558 ^ w7495;
	assign w48920 = w45640 ^ w7310;
	assign w47372 = w48920 ^ w1572;
	assign w33758 = w47372 ^ w47366;
	assign w33835 = w33752 ^ w33758;
	assign w33838 = w47367 ^ w33758;
	assign w7435 = w7558 ^ w7496;
	assign w7426 = w7558 ^ w7536;
	assign w7425 = w7426 ^ w7427;
	assign w48928 = w45268 ^ w7435;
	assign w48913 = ~w7425;
	assign w47380 = w48912 ^ w1564;
	assign w19286 = w47380 ^ w47374;
	assign w19366 = w47375 ^ w19286;
	assign w19365 = w47380 ^ w19241;
	assign w19351 = w47380 & w19365;
	assign w47364 = w48928 ^ w1580;
	assign w19152 = w47364 ^ w47358;
	assign w19222 = w19152 ^ w19147;
	assign w19232 = w47359 ^ w19152;
	assign w19228 = w47363 ^ w19232;
	assign w19231 = w47364 ^ w19107;
	assign w19217 = w47364 & w19231;
	assign w19215 = w19232 & w19228;
	assign w47355 = w48937 ^ w1589;
	assign w31288 = w47355 ^ w31292;
	assign w31222 = w47355 ^ w47354;
	assign w31287 = w31222 ^ w31289;
	assign w31295 = w47349 ^ w47355;
	assign w31275 = w31292 & w31288;
	assign w47379 = w48913 ^ w1565;
	assign w19279 = w47379 ^ w47377;
	assign w19281 = w47378 ^ w19279;
	assign w19357 = w47374 ^ w19281;
	assign w19354 = w47375 ^ w19281;
	assign w19356 = w19286 ^ w19281;
	assign w19362 = w47379 ^ w19366;
	assign w19296 = w47379 ^ w47378;
	assign w19349 = w19366 & w19362;
	assign w45912 = ~w7148;
	assign w7046 = w45912 ^ w48860;
	assign w48754 = w7045 ^ w7046;
	assign w7043 = w45912 ^ w48861;
	assign w47465 = w48754 ^ w1416;
	assign w34130 = w47465 ^ w47466;
	assign w48755 = w7042 ^ w7043;
	assign w47464 = w48755 ^ w1417;
	assign w34156 = w47464 ^ w47462;
	assign w34242 = w47464 ^ w47461;
	assign w34244 = w47466 ^ w47464;
	assign w34229 = w34154 ^ w34244;
	assign w34116 = w34156 ^ w34154;
	assign w34115 = w34156 ^ w47463;
	assign w34239 = w47468 ^ w34115;
	assign w34225 = w47468 & w34239;
	assign w34220 = w34244 & w34229;
	assign w7050 = w45912 ^ w45456;
	assign w7048 = w7049 ^ w7050;
	assign w48752 = ~w7048;
	assign w47467 = w48752 ^ w1414;
	assign w34153 = w47467 ^ w47465;
	assign w34155 = w47466 ^ w34153;
	assign w34231 = w47462 ^ w34155;
	assign w34228 = w47463 ^ w34155;
	assign w34230 = w34160 ^ w34155;
	assign w34236 = w47467 ^ w34240;
	assign w34234 = w34153 ^ w34242;
	assign w34233 = w47468 ^ w34234;
	assign w34170 = w47467 ^ w47466;
	assign w34235 = w34170 ^ w34237;
	assign w34238 = w34242 ^ w34170;
	assign w34232 = w34153 ^ w34116;
	assign w34243 = w47461 ^ w47467;
	assign w34227 = w34234 & w34238;
	assign w34159 = w34227 ^ w34156;
	assign w34226 = w34235 & w34233;
	assign w34177 = w34220 ^ w34226;
	assign w34224 = w34243 & w34228;
	assign w34158 = w34224 ^ w34154;
	assign w34223 = w34240 & w34236;
	assign w34222 = w34237 & w34230;
	assign w34221 = w34242 & w34231;
	assign w34157 = w34221 ^ w34155;
	assign w34163 = w34159 ^ w34157;
	assign w34168 = w47461 ^ w34163;
	assign w34218 = w34177 ^ w34168;
	assign w34129 = w34220 ^ w34221;
	assign w34176 = w34129 ^ w34130;
	assign w34175 = w34176 ^ w34158;
	assign w34217 = w34223 ^ w34175;
	assign w34219 = w34241 & w34232;
	assign w34214 = w34218 & w34217;
	assign w44800 = w34219 ^ w34225;
	assign w34169 = w44800 ^ w34154;
	assign w34215 = w34177 ^ w34169;
	assign w34131 = w34163 ^ w44800;
	assign w34174 = w47463 ^ w34131;
	assign w34209 = w34214 ^ w34174;
	assign w44801 = w34219 ^ w34222;
	assign w34172 = w34220 ^ w44801;
	assign w34128 = w34223 ^ w34172;
	assign w34210 = w47467 ^ w34128;
	assign w34208 = w34209 & w34210;
	assign w34127 = w34208 ^ w34172;
	assign w34126 = w34208 ^ w34225;
	assign w34121 = w34126 ^ w34222;
	assign w34206 = w34214 ^ w34208;
	assign w34132 = w34158 ^ w44801;
	assign w34216 = w34132 ^ w34157;
	assign w34207 = w34208 ^ w34216;
	assign w34213 = w34214 ^ w34216;
	assign w34212 = w34215 & w34213;
	assign w34211 = w34212 ^ w34174;
	assign w34123 = w34212 ^ w34224;
	assign w34119 = w34123 ^ w34159;
	assign w34122 = w47461 ^ w34119;
	assign w34199 = w34121 ^ w34122;
	assign w34120 = w34212 ^ w34168;
	assign w34118 = w47463 ^ w34119;
	assign w34205 = w34216 & w34206;
	assign w34203 = w34205 ^ w34213;
	assign w34202 = w34211 & w34203;
	assign w34167 = w34202 ^ w34177;
	assign w34201 = w34167 ^ w34169;
	assign w34125 = w34202 ^ w34226;
	assign w34198 = w34167 ^ w34120;
	assign w34193 = w34207 & w47468;
	assign w34192 = w34198 & w34228;
	assign w34191 = w34201 & w34240;
	assign w34190 = w34211 & w34230;
	assign w34134 = w34190 ^ w34191;
	assign w34189 = w34199 & w34231;
	assign w34184 = w34207 & w34239;
	assign w34183 = w34198 & w34243;
	assign w34150 = w34192 ^ w34183;
	assign w34182 = w34201 & w34236;
	assign w34152 = w34190 ^ w34182;
	assign w34181 = w34211 & w34237;
	assign w34180 = w34199 & w34242;
	assign w44802 = w34191 ^ w34192;
	assign w44804 = w34205 ^ w34223;
	assign w34164 = w47467 ^ w44804;
	assign w34204 = w34164 ^ w34127;
	assign w34185 = w34204 & w34235;
	assign w34194 = w34204 & w34233;
	assign w34117 = w34164 ^ w34125;
	assign w34124 = w34154 ^ w34117;
	assign w34200 = w34121 ^ w34124;
	assign w34187 = w34200 & w34232;
	assign w34165 = w34183 ^ w34187;
	assign w34143 = ~w34165;
	assign w34142 = w34143 ^ w34181;
	assign w34196 = w34117 ^ w34118;
	assign w34179 = w34196 & w34244;
	assign w34178 = w34200 & w34241;
	assign w34144 = w34189 ^ w34178;
	assign w34140 = ~w34144;
	assign w43595 = w34179 ^ w34180;
	assign w34161 = w34185 ^ w43595;
	assign w34148 = w34152 ^ w43595;
	assign w34147 = w34143 ^ w34148;
	assign w34188 = w34196 & w34229;
	assign w34145 = w34188 ^ w34189;
	assign w34173 = w34188 ^ w44802;
	assign w34139 = w34184 ^ w34173;
	assign w34136 = ~w34139;
	assign w34133 = w34189 ^ w34173;
	assign w34149 = w34188 ^ w34191;
	assign w34146 = ~w34149;
	assign w34247 = w34146 ^ w34147;
	assign w34197 = w44804 ^ w34175;
	assign w34195 = w34197 & w34234;
	assign w34186 = w34197 & w34238;
	assign w34162 = w34186 ^ w34161;
	assign w34166 = w34194 ^ w34162;
	assign w34171 = w34195 ^ w34166;
	assign w49103 = w44802 ^ w34171;
	assign w34246 = w34171 ^ w34145;
	assign w34135 = w34193 ^ w34166;
	assign w49102 = w34134 ^ w34135;
	assign w49104 = w34162 ^ w34133;
	assign w7503 = w49104 ^ w49108;
	assign w7242 = w7503 ^ w49105;
	assign w7240 = w7503 ^ w45723;
	assign w7508 = w49102 ^ w49106;
	assign w49011 = w7576 ^ w7508;
	assign w47281 = w49011 ^ w1472;
	assign w7489 = w49100 ^ w49104;
	assign w7480 = w49104 ^ w20042;
	assign w7478 = w7538 ^ w7489;
	assign w49016 = w45443 ^ w7478;
	assign w7486 = w7500 ^ w49103;
	assign w49012 = w7485 ^ w7486;
	assign w47280 = w49012 ^ w1473;
	assign w7442 = w7511 ^ w7489;
	assign w49039 = w49108 ^ w7442;
	assign w47253 = w49039 ^ w1499;
	assign w7460 = w7503 ^ w49111;
	assign w7454 = w7489 ^ w49112;
	assign w7447 = w7508 ^ w7506;
	assign w7293 = w49102 ^ w7294;
	assign w47276 = w49016 ^ w1477;
	assign w44803 = w34193 ^ w34195;
	assign w34151 = w44803 ^ w34148;
	assign w34248 = w34150 ^ w34151;
	assign w34138 = w34142 ^ w44803;
	assign w34141 = w34180 ^ w34138;
	assign w34245 = w34140 ^ w34141;
	assign w34137 = w34161 ^ w34138;
	assign w49101 = w34136 ^ w34137;
	assign w7243 = w49102 ^ w49101;
	assign w7582 = w7242 ^ w7243;
	assign w49027 = w7582 ^ w7514;
	assign w7528 = w49096 ^ w49101;
	assign w7473 = w7528 ^ w7514;
	assign w7471 = ~w7473;
	assign w7461 = w7528 ^ w49109;
	assign w7298 = w45723 ^ w49101;
	assign w49010 = w7297 ^ w7298;
	assign w47282 = w49010 ^ w1471;
	assign w18834 = w47282 ^ w47280;
	assign w18720 = w47281 ^ w47282;
	assign w7449 = w7528 ^ w7518;
	assign w49034 = w49105 ^ w7449;
	assign w47258 = w49034 ^ w1494;
	assign w7711 = w47253 ^ w47258;
	assign w47265 = w49027 ^ w1488;
	assign w7554 = w49098 ^ w49103;
	assign w49036 = w7560 ^ w7554;
	assign w47256 = w49036 ^ w1496;
	assign w7712 = w47256 ^ w47253;
	assign w7714 = w47258 ^ w47256;
	assign w7470 = w7554 ^ w7523;
	assign w49021 = w45436 ^ w7470;
	assign w47271 = w49021 ^ w1482;
	assign w7459 = w7554 ^ w7508;
	assign w49028 = w7459 ^ w7460;
	assign w47264 = w49028 ^ w1489;
	assign w45786 = ~w34245;
	assign w7513 = w45786 ^ w45436;
	assign w7466 = w7511 ^ w45786;
	assign w7465 = w7466 ^ w7467;
	assign w49022 = ~w7465;
	assign w7484 = ~w7513;
	assign w7482 = w7484 ^ w45729;
	assign w49013 = w7482 ^ w7483;
	assign w47279 = w49013 ^ w1474;
	assign w7445 = w7513 ^ w7505;
	assign w49037 = w45449 ^ w7445;
	assign w7458 = w45786 ^ w49103;
	assign w49029 = w7457 ^ w7458;
	assign w47263 = w49029 ^ w1490;
	assign w47255 = w49037 ^ w1497;
	assign w7624 = w47255 ^ w47253;
	assign w7699 = w7624 ^ w7714;
	assign w47270 = w49022 ^ w1483;
	assign w34026 = w47276 ^ w47270;
	assign w34106 = w47271 ^ w34026;
	assign w7690 = w7714 & w7699;
	assign w45787 = ~w34246;
	assign w49014 = w45787 ^ w7481;
	assign w47278 = w49014 ^ w1475;
	assign w18746 = w47280 ^ w47278;
	assign w18705 = w18746 ^ w47279;
	assign w7553 = w49099 ^ w45787;
	assign w7464 = w7553 ^ w7488;
	assign w49023 = w49100 ^ w7464;
	assign w7443 = w7553 ^ w45729;
	assign w7456 = w7553 ^ w7513;
	assign w49030 = w45722 ^ w7456;
	assign w47262 = w49030 ^ w1491;
	assign w18612 = w47264 ^ w47262;
	assign w18571 = w18612 ^ w47263;
	assign w49038 = w7443 ^ w7444;
	assign w47254 = w49038 ^ w1498;
	assign w7626 = w47256 ^ w47254;
	assign w7585 = w7626 ^ w47255;
	assign w7586 = w7626 ^ w7624;
	assign w47269 = w49023 ^ w1484;
	assign w34020 = w47271 ^ w47269;
	assign w34103 = w34020 ^ w34026;
	assign w7455 = w45437 ^ w45787;
	assign w49031 = w7454 ^ w7455;
	assign w47261 = w49031 ^ w1492;
	assign w18610 = w47263 ^ w47261;
	assign w18698 = w47264 ^ w47261;
	assign w18572 = w18612 ^ w18610;
	assign w45788 = ~w34247;
	assign w7255 = w45724 ^ w45788;
	assign w7577 = w7254 ^ w7255;
	assign w49009 = w7577 ^ w7518;
	assign w47283 = w49009 ^ w1470;
	assign w18743 = w47283 ^ w47281;
	assign w18745 = w47282 ^ w18743;
	assign w18821 = w47278 ^ w18745;
	assign w18818 = w47279 ^ w18745;
	assign w18760 = w47283 ^ w47282;
	assign w7543 = w45442 ^ w45788;
	assign w7474 = w7543 ^ w7506;
	assign w49018 = w49096 ^ w7474;
	assign w7462 = w45430 ^ w45788;
	assign w49026 = w7461 ^ w7462;
	assign w7452 = ~w7543;
	assign w7450 = w7452 ^ w7538;
	assign w47266 = w49026 ^ w1487;
	assign w18700 = w47266 ^ w47264;
	assign w18685 = w18610 ^ w18700;
	assign w18586 = w47265 ^ w47266;
	assign w18697 = w47261 ^ w47266;
	assign w18676 = w18700 & w18685;
	assign w47274 = w49018 ^ w1479;
	assign w34107 = w47269 ^ w47274;
	assign w45789 = ~w34248;
	assign w7241 = w45431 ^ w45789;
	assign w7583 = w7240 ^ w7241;
	assign w49025 = w7583 ^ w7543;
	assign w7551 = w45443 ^ w45789;
	assign w7463 = w7551 ^ w7503;
	assign w49024 = w45724 ^ w7463;
	assign w7476 = w7551 ^ w7518;
	assign w49008 = w45789 ^ w7299;
	assign w47284 = w49008 ^ w1469;
	assign w18750 = w47284 ^ w47278;
	assign w18820 = w18750 ^ w18745;
	assign w18830 = w47279 ^ w18750;
	assign w18826 = w47283 ^ w18830;
	assign w18829 = w47284 ^ w18705;
	assign w18815 = w47284 & w18829;
	assign w18813 = w18830 & w18826;
	assign w7453 = w7551 ^ w7488;
	assign w49032 = w45431 ^ w7453;
	assign w47260 = w49032 ^ w1493;
	assign w7709 = w47260 ^ w7585;
	assign w7695 = w47260 & w7709;
	assign w7630 = w47260 ^ w47254;
	assign w7710 = w47255 ^ w7630;
	assign w7707 = w7624 ^ w7630;
	assign w47267 = w49025 ^ w1486;
	assign w18609 = w47267 ^ w47265;
	assign w18611 = w47266 ^ w18609;
	assign w18687 = w47262 ^ w18611;
	assign w18684 = w47263 ^ w18611;
	assign w18690 = w18609 ^ w18698;
	assign w18626 = w47267 ^ w47266;
	assign w18694 = w18698 ^ w18626;
	assign w18688 = w18609 ^ w18572;
	assign w18699 = w47261 ^ w47267;
	assign w18683 = w18690 & w18694;
	assign w18615 = w18683 ^ w18612;
	assign w18680 = w18699 & w18684;
	assign w18614 = w18680 ^ w18610;
	assign w18677 = w18698 & w18687;
	assign w18613 = w18677 ^ w18611;
	assign w18619 = w18615 ^ w18613;
	assign w18624 = w47261 ^ w18619;
	assign w18585 = w18676 ^ w18677;
	assign w18632 = w18585 ^ w18586;
	assign w18631 = w18632 ^ w18614;
	assign w18675 = w18697 & w18688;
	assign w47268 = w49024 ^ w1485;
	assign w18689 = w47268 ^ w18690;
	assign w18616 = w47268 ^ w47262;
	assign w18686 = w18616 ^ w18611;
	assign w18693 = w18610 ^ w18616;
	assign w18691 = w18626 ^ w18693;
	assign w18696 = w47263 ^ w18616;
	assign w18692 = w47267 ^ w18696;
	assign w18695 = w47268 ^ w18571;
	assign w18682 = w18691 & w18689;
	assign w18633 = w18676 ^ w18682;
	assign w18674 = w18633 ^ w18624;
	assign w18681 = w47268 & w18695;
	assign w18679 = w18696 & w18692;
	assign w18673 = w18679 ^ w18631;
	assign w18678 = w18693 & w18686;
	assign w18670 = w18674 & w18673;
	assign w44148 = w18675 ^ w18678;
	assign w18588 = w18614 ^ w44148;
	assign w18672 = w18588 ^ w18613;
	assign w18669 = w18670 ^ w18672;
	assign w18628 = w18676 ^ w44148;
	assign w18584 = w18679 ^ w18628;
	assign w18666 = w47267 ^ w18584;
	assign w44151 = w18675 ^ w18681;
	assign w18587 = w18619 ^ w44151;
	assign w18630 = w47263 ^ w18587;
	assign w18665 = w18670 ^ w18630;
	assign w18664 = w18665 & w18666;
	assign w18662 = w18670 ^ w18664;
	assign w18583 = w18664 ^ w18628;
	assign w18582 = w18664 ^ w18681;
	assign w18577 = w18582 ^ w18678;
	assign w18661 = w18672 & w18662;
	assign w18659 = w18661 ^ w18669;
	assign w44150 = w18661 ^ w18679;
	assign w18653 = w44150 ^ w18631;
	assign w18642 = w18653 & w18694;
	assign w18651 = w18653 & w18690;
	assign w18620 = w47267 ^ w44150;
	assign w18660 = w18620 ^ w18583;
	assign w18650 = w18660 & w18689;
	assign w18641 = w18660 & w18691;
	assign w18663 = w18664 ^ w18672;
	assign w18649 = w18663 & w47268;
	assign w18640 = w18663 & w18695;
	assign w18625 = w44151 ^ w18610;
	assign w18671 = w18633 ^ w18625;
	assign w18668 = w18671 & w18669;
	assign w18667 = w18668 ^ w18630;
	assign w18579 = w18668 ^ w18680;
	assign w18575 = w18579 ^ w18615;
	assign w18578 = w47261 ^ w18575;
	assign w18655 = w18577 ^ w18578;
	assign w18576 = w18668 ^ w18624;
	assign w18574 = w47263 ^ w18575;
	assign w18658 = w18667 & w18659;
	assign w18623 = w18658 ^ w18633;
	assign w18657 = w18623 ^ w18625;
	assign w18581 = w18658 ^ w18682;
	assign w18573 = w18620 ^ w18581;
	assign w18580 = w18610 ^ w18573;
	assign w18656 = w18577 ^ w18580;
	assign w18654 = w18623 ^ w18576;
	assign w18652 = w18573 ^ w18574;
	assign w18648 = w18654 & w18684;
	assign w18647 = w18657 & w18696;
	assign w18646 = w18667 & w18686;
	assign w18590 = w18646 ^ w18647;
	assign w18645 = w18655 & w18687;
	assign w18644 = w18652 & w18685;
	assign w18605 = w18644 ^ w18647;
	assign w18602 = ~w18605;
	assign w18601 = w18644 ^ w18645;
	assign w18643 = w18656 & w18688;
	assign w18639 = w18654 & w18699;
	assign w18621 = w18639 ^ w18643;
	assign w18606 = w18648 ^ w18639;
	assign w18599 = ~w18621;
	assign w18638 = w18657 & w18692;
	assign w18608 = w18646 ^ w18638;
	assign w18637 = w18667 & w18693;
	assign w18598 = w18599 ^ w18637;
	assign w18636 = w18655 & w18698;
	assign w18635 = w18652 & w18700;
	assign w18634 = w18656 & w18697;
	assign w18600 = w18645 ^ w18634;
	assign w18596 = ~w18600;
	assign w44149 = w18635 ^ w18636;
	assign w18617 = w18641 ^ w44149;
	assign w18618 = w18642 ^ w18617;
	assign w18622 = w18650 ^ w18618;
	assign w18591 = w18649 ^ w18622;
	assign w49253 = w18590 ^ w18591;
	assign w18627 = w18651 ^ w18622;
	assign w18702 = w18627 ^ w18601;
	assign w18604 = w18608 ^ w44149;
	assign w18603 = w18599 ^ w18604;
	assign w18703 = w18602 ^ w18603;
	assign w49251 = ~w18703;
	assign w44152 = w18647 ^ w18648;
	assign w49254 = w44152 ^ w18627;
	assign w18629 = w18644 ^ w44152;
	assign w18595 = w18640 ^ w18629;
	assign w18592 = ~w18595;
	assign w18589 = w18645 ^ w18629;
	assign w49255 = w18618 ^ w18589;
	assign w44153 = w18649 ^ w18651;
	assign w18607 = w44153 ^ w18604;
	assign w18704 = w18606 ^ w18607;
	assign w18594 = w18598 ^ w44153;
	assign w18597 = w18636 ^ w18594;
	assign w18701 = w18596 ^ w18597;
	assign w18593 = w18617 ^ w18594;
	assign w49252 = w18592 ^ w18593;
	assign w7770 = ~w49252;
	assign w7769 = w49253 ^ w7770;
	assign w45407 = ~w18701;
	assign w45408 = ~w18702;
	assign w45409 = ~w18704;
	assign w45913 = ~w7146;
	assign w6960 = w45913 ^ w48889;
	assign w6963 = w45913 ^ w48888;
	assign w48802 = w6962 ^ w6963;
	assign w6968 = w45913 ^ w45555;
	assign w48800 = w6967 ^ w6968;
	assign w48803 = w6959 ^ w6960;
	assign w47416 = w48803 ^ w1401;
	assign w28394 = w47416 ^ w47414;
	assign w28480 = w47416 ^ w47413;
	assign w28482 = w47418 ^ w47416;
	assign w28467 = w28392 ^ w28482;
	assign w28354 = w28394 ^ w28392;
	assign w28353 = w28394 ^ w47415;
	assign w28477 = w47420 ^ w28353;
	assign w28463 = w47420 & w28477;
	assign w28458 = w28482 & w28467;
	assign w47417 = w48802 ^ w1400;
	assign w28368 = w47417 ^ w47418;
	assign w47419 = w48800 ^ w1398;
	assign w28391 = w47419 ^ w47417;
	assign w28393 = w47418 ^ w28391;
	assign w28469 = w47414 ^ w28393;
	assign w28466 = w47415 ^ w28393;
	assign w28468 = w28398 ^ w28393;
	assign w28474 = w47419 ^ w28478;
	assign w28472 = w28391 ^ w28480;
	assign w28471 = w47420 ^ w28472;
	assign w28408 = w47419 ^ w47418;
	assign w28473 = w28408 ^ w28475;
	assign w28476 = w28480 ^ w28408;
	assign w28470 = w28391 ^ w28354;
	assign w28481 = w47413 ^ w47419;
	assign w28465 = w28472 & w28476;
	assign w28397 = w28465 ^ w28394;
	assign w28464 = w28473 & w28471;
	assign w28415 = w28458 ^ w28464;
	assign w28462 = w28481 & w28466;
	assign w28396 = w28462 ^ w28392;
	assign w28461 = w28478 & w28474;
	assign w28460 = w28475 & w28468;
	assign w28459 = w28480 & w28469;
	assign w28395 = w28459 ^ w28393;
	assign w28401 = w28397 ^ w28395;
	assign w28406 = w47413 ^ w28401;
	assign w28456 = w28415 ^ w28406;
	assign w28367 = w28458 ^ w28459;
	assign w28414 = w28367 ^ w28368;
	assign w28413 = w28414 ^ w28396;
	assign w28455 = w28461 ^ w28413;
	assign w28457 = w28479 & w28470;
	assign w28452 = w28456 & w28455;
	assign w44557 = w28457 ^ w28463;
	assign w28369 = w28401 ^ w44557;
	assign w28412 = w47415 ^ w28369;
	assign w28447 = w28452 ^ w28412;
	assign w28407 = w44557 ^ w28392;
	assign w28453 = w28415 ^ w28407;
	assign w44558 = w28457 ^ w28460;
	assign w28410 = w28458 ^ w44558;
	assign w28366 = w28461 ^ w28410;
	assign w28448 = w47419 ^ w28366;
	assign w28446 = w28447 & w28448;
	assign w28365 = w28446 ^ w28410;
	assign w28444 = w28452 ^ w28446;
	assign w28364 = w28446 ^ w28463;
	assign w28359 = w28364 ^ w28460;
	assign w28370 = w28396 ^ w44558;
	assign w28454 = w28370 ^ w28395;
	assign w28445 = w28446 ^ w28454;
	assign w28451 = w28452 ^ w28454;
	assign w28450 = w28453 & w28451;
	assign w28449 = w28450 ^ w28412;
	assign w28361 = w28450 ^ w28462;
	assign w28357 = w28361 ^ w28397;
	assign w28360 = w47413 ^ w28357;
	assign w28437 = w28359 ^ w28360;
	assign w28358 = w28450 ^ w28406;
	assign w28356 = w47415 ^ w28357;
	assign w28443 = w28454 & w28444;
	assign w28441 = w28443 ^ w28451;
	assign w28440 = w28449 & w28441;
	assign w28405 = w28440 ^ w28415;
	assign w28439 = w28405 ^ w28407;
	assign w28363 = w28440 ^ w28464;
	assign w28436 = w28405 ^ w28358;
	assign w28431 = w28445 & w47420;
	assign w28430 = w28436 & w28466;
	assign w28429 = w28439 & w28478;
	assign w28428 = w28449 & w28468;
	assign w28372 = w28428 ^ w28429;
	assign w28427 = w28437 & w28469;
	assign w28422 = w28445 & w28477;
	assign w28421 = w28436 & w28481;
	assign w28388 = w28430 ^ w28421;
	assign w28420 = w28439 & w28474;
	assign w28390 = w28428 ^ w28420;
	assign w28419 = w28449 & w28475;
	assign w28418 = w28437 & w28480;
	assign w44560 = w28429 ^ w28430;
	assign w44562 = w28443 ^ w28461;
	assign w28435 = w44562 ^ w28413;
	assign w28433 = w28435 & w28472;
	assign w44561 = w28431 ^ w28433;
	assign w28424 = w28435 & w28476;
	assign w28402 = w47419 ^ w44562;
	assign w28442 = w28402 ^ w28365;
	assign w28355 = w28402 ^ w28363;
	assign w28362 = w28392 ^ w28355;
	assign w28438 = w28359 ^ w28362;
	assign w28434 = w28355 ^ w28356;
	assign w28432 = w28442 & w28471;
	assign w28426 = w28434 & w28467;
	assign w28411 = w28426 ^ w44560;
	assign w28387 = w28426 ^ w28429;
	assign w28384 = ~w28387;
	assign w28383 = w28426 ^ w28427;
	assign w28377 = w28422 ^ w28411;
	assign w28374 = ~w28377;
	assign w28371 = w28427 ^ w28411;
	assign w28425 = w28438 & w28470;
	assign w28403 = w28421 ^ w28425;
	assign w28381 = ~w28403;
	assign w28380 = w28381 ^ w28419;
	assign w28376 = w28380 ^ w44561;
	assign w28379 = w28418 ^ w28376;
	assign w28423 = w28442 & w28473;
	assign w28417 = w28434 & w28482;
	assign w28416 = w28438 & w28479;
	assign w28382 = w28427 ^ w28416;
	assign w28378 = ~w28382;
	assign w28483 = w28378 ^ w28379;
	assign w44559 = w28417 ^ w28418;
	assign w28399 = w28423 ^ w44559;
	assign w28375 = w28399 ^ w28376;
	assign w49092 = w28374 ^ w28375;
	assign w28400 = w28424 ^ w28399;
	assign w49095 = w28400 ^ w28371;
	assign w28404 = w28432 ^ w28400;
	assign w28373 = w28431 ^ w28404;
	assign w49093 = w28372 ^ w28373;
	assign w28409 = w28433 ^ w28404;
	assign w28484 = w28409 ^ w28383;
	assign w7490 = w49091 ^ w49095;
	assign w7498 = w49080 ^ w49095;
	assign w7271 = w7498 ^ w49093;
	assign w7267 = ~w7498;
	assign w7268 = w7267 ^ w49092;
	assign w7530 = w49089 ^ w49093;
	assign w7540 = w49088 ^ w49092;
	assign w7353 = ~w7540;
	assign w49094 = w44560 ^ w28409;
	assign w7521 = w49090 ^ w49094;
	assign w28386 = w28390 ^ w44559;
	assign w28389 = w44561 ^ w28386;
	assign w28486 = w28388 ^ w28389;
	assign w28385 = w28381 ^ w28386;
	assign w28485 = w28384 ^ w28385;
	assign w45642 = ~w28483;
	assign w7515 = w45440 ^ w45642;
	assign w7350 = w7515 ^ w49094;
	assign w7348 = ~w7350;
	assign w45643 = ~w28484;
	assign w7340 = w7490 ^ w45643;
	assign w7504 = w45441 ^ w45643;
	assign w7343 = w7504 ^ w45642;
	assign w45644 = ~w28485;
	assign w7351 = w7353 ^ w45644;
	assign w7544 = w45434 ^ w45644;
	assign w45645 = ~w28486;
	assign w7265 = w7267 ^ w45645;
	assign w7552 = w45435 ^ w45645;
	assign w7354 = w7552 ^ w7498;
	assign w45914 = ~w7145;
	assign w6948 = w45914 ^ w48896;
	assign w7217 = w6948 ^ w6949;
	assign w48819 = w7217 ^ w7161;
	assign w47400 = w48819 ^ w2022;
	assign w13340 = w47402 ^ w47400;
	assign w13325 = w13250 ^ w13340;
	assign w13316 = w13340 & w13325;
	assign w13338 = w47400 ^ w47397;
	assign w7128 = w45914 ^ w48905;
	assign w7133 = w45914 ^ w45559;
	assign w7131 = w7132 ^ w7133;
	assign w48816 = ~w7131;
	assign w47403 = w48816 ^ w2019;
	assign w13332 = w47403 ^ w13336;
	assign w13266 = w47403 ^ w47402;
	assign w13331 = w13266 ^ w13333;
	assign w13339 = w47397 ^ w47403;
	assign w13319 = w13336 & w13332;
	assign w13334 = w13338 ^ w13266;
	assign w48818 = w7127 ^ w7128;
	assign w47401 = w48818 ^ w2021;
	assign w13226 = w47401 ^ w47402;
	assign w13249 = w47403 ^ w47401;
	assign w13330 = w13249 ^ w13338;
	assign w13323 = w13330 & w13334;
	assign w13329 = w47404 ^ w13330;
	assign w13322 = w13331 & w13329;
	assign w13273 = w13316 ^ w13322;
	assign w13251 = w47402 ^ w13249;
	assign w13324 = w47399 ^ w13251;
	assign w13327 = w47398 ^ w13251;
	assign w13326 = w13256 ^ w13251;
	assign w13320 = w13339 & w13324;
	assign w13318 = w13333 & w13326;
	assign w13317 = w13338 & w13327;
	assign w13225 = w13316 ^ w13317;
	assign w13272 = w13225 ^ w13226;
	assign w13253 = w13317 ^ w13251;
	assign w13252 = w47400 ^ w47398;
	assign w13255 = w13323 ^ w13252;
	assign w13259 = w13255 ^ w13253;
	assign w13211 = w13252 ^ w47399;
	assign w13335 = w47404 ^ w13211;
	assign w13321 = w47404 & w13335;
	assign w13212 = w13252 ^ w13250;
	assign w13328 = w13249 ^ w13212;
	assign w13315 = w13337 & w13328;
	assign w13264 = w47397 ^ w13259;
	assign w13314 = w13273 ^ w13264;
	assign w43926 = w13315 ^ w13321;
	assign w13265 = w43926 ^ w13250;
	assign w13311 = w13273 ^ w13265;
	assign w13227 = w13259 ^ w43926;
	assign w13270 = w47399 ^ w13227;
	assign w43927 = w13315 ^ w13318;
	assign w13268 = w13316 ^ w43927;
	assign w13224 = w13319 ^ w13268;
	assign w13306 = w47403 ^ w13224;
	assign w13254 = w13320 ^ w13250;
	assign w13228 = w13254 ^ w43927;
	assign w13312 = w13228 ^ w13253;
	assign w13271 = w13272 ^ w13254;
	assign w13313 = w13319 ^ w13271;
	assign w13310 = w13314 & w13313;
	assign w13309 = w13310 ^ w13312;
	assign w13308 = w13311 & w13309;
	assign w13219 = w13308 ^ w13320;
	assign w13215 = w13219 ^ w13255;
	assign w13218 = w47397 ^ w13215;
	assign w13216 = w13308 ^ w13264;
	assign w13214 = w47399 ^ w13215;
	assign w13307 = w13308 ^ w13270;
	assign w13286 = w13307 & w13326;
	assign w13277 = w13307 & w13333;
	assign w13305 = w13310 ^ w13270;
	assign w13304 = w13305 & w13306;
	assign w13303 = w13304 ^ w13312;
	assign w13223 = w13304 ^ w13268;
	assign w13222 = w13304 ^ w13321;
	assign w13302 = w13310 ^ w13304;
	assign w13289 = w13303 & w47404;
	assign w13280 = w13303 & w13335;
	assign w13301 = w13312 & w13302;
	assign w13299 = w13301 ^ w13309;
	assign w13298 = w13307 & w13299;
	assign w13221 = w13298 ^ w13322;
	assign w13217 = w13222 ^ w13318;
	assign w13295 = w13217 ^ w13218;
	assign w13285 = w13295 & w13327;
	assign w13276 = w13295 & w13338;
	assign w13263 = w13298 ^ w13273;
	assign w13294 = w13263 ^ w13216;
	assign w13297 = w13263 ^ w13265;
	assign w13279 = w13294 & w13339;
	assign w13288 = w13294 & w13324;
	assign w13287 = w13297 & w13336;
	assign w13230 = w13286 ^ w13287;
	assign w13278 = w13297 & w13332;
	assign w13246 = w13288 ^ w13279;
	assign w13248 = w13286 ^ w13278;
	assign w43928 = w13287 ^ w13288;
	assign w43930 = w13301 ^ w13319;
	assign w13260 = w47403 ^ w43930;
	assign w13300 = w13260 ^ w13223;
	assign w13290 = w13300 & w13329;
	assign w13281 = w13300 & w13331;
	assign w13213 = w13260 ^ w13221;
	assign w13220 = w13250 ^ w13213;
	assign w13296 = w13217 ^ w13220;
	assign w13283 = w13296 & w13328;
	assign w13274 = w13296 & w13337;
	assign w13240 = w13285 ^ w13274;
	assign w13261 = w13279 ^ w13283;
	assign w13239 = ~w13261;
	assign w13238 = w13239 ^ w13277;
	assign w13236 = ~w13240;
	assign w13292 = w13213 ^ w13214;
	assign w13284 = w13292 & w13325;
	assign w13245 = w13284 ^ w13287;
	assign w13242 = ~w13245;
	assign w13241 = w13284 ^ w13285;
	assign w13275 = w13292 & w13340;
	assign w43533 = w13275 ^ w13276;
	assign w13257 = w13281 ^ w43533;
	assign w13244 = w13248 ^ w43533;
	assign w13243 = w13239 ^ w13244;
	assign w13343 = w13242 ^ w13243;
	assign w49064 = ~w13343;
	assign w7531 = w45547 ^ w49064;
	assign w7247 = w13343 ^ w45548;
	assign w7580 = w7246 ^ w7247;
	assign w13293 = w43930 ^ w13271;
	assign w13291 = w13293 & w13330;
	assign w13282 = w13293 & w13334;
	assign w13258 = w13282 ^ w13257;
	assign w13262 = w13290 ^ w13258;
	assign w13231 = w13289 ^ w13262;
	assign w49066 = w13230 ^ w13231;
	assign w13267 = w13291 ^ w13262;
	assign w13342 = w13267 ^ w13241;
	assign w7251 = ~w49066;
	assign w7250 = w7251 ^ w49060;
	assign w7579 = w7249 ^ w7250;
	assign w7524 = w49061 ^ w49066;
	assign w7388 = ~w7524;
	assign w49067 = w43928 ^ w13267;
	assign w7253 = w49067 ^ w49061;
	assign w7578 = w7252 ^ w7253;
	assign w7520 = w49062 ^ w49067;
	assign w7362 = ~w7520;
	assign w43929 = w13289 ^ w13291;
	assign w13247 = w43929 ^ w13244;
	assign w13344 = w13246 ^ w13247;
	assign w13234 = w13238 ^ w43929;
	assign w13237 = w13276 ^ w13234;
	assign w13341 = w13236 ^ w13237;
	assign w13233 = w13257 ^ w13234;
	assign w45262 = ~w13342;
	assign w45263 = ~w13344;
	assign w7532 = w45548 ^ w45263;
	assign w45269 = ~w13341;
	assign w7374 = w45262 ^ w45269;
	assign w7516 = w45553 ^ w45269;
	assign w7377 = w7516 ^ w45733;
	assign w7384 = w7516 ^ w7510;
	assign w7375 = ~w7377;
	assign w7404 = w45269 ^ w49062;
	assign w13269 = w13284 ^ w43928;
	assign w13235 = w13280 ^ w13269;
	assign w13229 = w13285 ^ w13269;
	assign w49068 = w13258 ^ w13229;
	assign w13232 = ~w13235;
	assign w49065 = w13232 ^ w13233;
	assign w7492 = w49063 ^ w49068;
	assign w7584 = ~w7492;
	assign w7390 = w7584 ^ w49061;
	assign w7394 = w7584 ^ w45547;
	assign w7527 = w49060 ^ w49065;
	assign w7380 = ~w7527;
	assign w7378 = w7380 ^ w49073;
	assign w7406 = w49065 ^ w45547;
	assign w7387 = w7584 ^ w49062;
	assign w7355 = w7492 ^ w45726;
	assign w45915 = ~w7151;
	assign w6939 = w45915 ^ w45793;
	assign w7221 = w6939 ^ w6940;
	assign w48720 = w7221 ^ w7213;
	assign w47499 = w48720 ^ w1446;
	assign w13600 = w47499 ^ w13604;
	assign w13517 = w47499 ^ w47497;
	assign w13519 = w47498 ^ w13517;
	assign w13594 = w13524 ^ w13519;
	assign w13534 = w47499 ^ w47498;
	assign w13599 = w13534 ^ w13601;
	assign w13587 = w13604 & w13600;
	assign w13586 = w13601 & w13594;
	assign w13607 = w47493 ^ w47499;
	assign w13595 = w47494 ^ w13519;
	assign w13592 = w47495 ^ w13519;
	assign w13588 = w13607 & w13592;
	assign w13522 = w13588 ^ w13518;
	assign w7096 = w45915 ^ w48841;
	assign w48723 = w7095 ^ w7096;
	assign w47496 = w48723 ^ w1449;
	assign w13608 = w47498 ^ w47496;
	assign w13520 = w47496 ^ w47494;
	assign w13593 = w13518 ^ w13608;
	assign w13606 = w47496 ^ w47493;
	assign w13602 = w13606 ^ w13534;
	assign w13598 = w13517 ^ w13606;
	assign w13597 = w47500 ^ w13598;
	assign w13585 = w13606 & w13595;
	assign w13521 = w13585 ^ w13519;
	assign w13479 = w13520 ^ w47495;
	assign w13480 = w13520 ^ w13518;
	assign w13603 = w47500 ^ w13479;
	assign w13591 = w13598 & w13602;
	assign w13523 = w13591 ^ w13520;
	assign w13527 = w13523 ^ w13521;
	assign w13532 = w47493 ^ w13527;
	assign w13590 = w13599 & w13597;
	assign w13589 = w47500 & w13603;
	assign w13596 = w13517 ^ w13480;
	assign w13583 = w13605 & w13596;
	assign w13584 = w13608 & w13593;
	assign w13493 = w13584 ^ w13585;
	assign w13540 = w13493 ^ w13494;
	assign w13541 = w13584 ^ w13590;
	assign w13582 = w13541 ^ w13532;
	assign w13539 = w13540 ^ w13522;
	assign w7075 = w45915 ^ w48858;
	assign w48734 = w7075 ^ w7076;
	assign w47485 = w48734 ^ w1460;
	assign w25176 = w47487 ^ w47485;
	assign w25251 = w25176 ^ w25266;
	assign w25264 = w47488 ^ w47485;
	assign w25260 = w25264 ^ w25192;
	assign w25259 = w25176 ^ w25182;
	assign w25257 = w25192 ^ w25259;
	assign w25256 = w25175 ^ w25264;
	assign w25255 = w47492 ^ w25256;
	assign w25138 = w25178 ^ w25176;
	assign w25254 = w25175 ^ w25138;
	assign w25265 = w47485 ^ w47491;
	assign w25263 = w47485 ^ w47490;
	assign w25249 = w25256 & w25260;
	assign w25181 = w25249 ^ w25178;
	assign w25248 = w25257 & w25255;
	assign w25246 = w25265 & w25250;
	assign w25180 = w25246 ^ w25176;
	assign w25244 = w25259 & w25252;
	assign w25243 = w25264 & w25253;
	assign w25179 = w25243 ^ w25177;
	assign w25185 = w25181 ^ w25179;
	assign w25190 = w47485 ^ w25185;
	assign w25242 = w25266 & w25251;
	assign w25199 = w25242 ^ w25248;
	assign w25240 = w25199 ^ w25190;
	assign w25151 = w25242 ^ w25243;
	assign w25198 = w25151 ^ w25152;
	assign w25197 = w25198 ^ w25180;
	assign w25239 = w25245 ^ w25197;
	assign w25241 = w25263 & w25254;
	assign w25236 = w25240 & w25239;
	assign w43937 = w13583 ^ w13589;
	assign w13533 = w43937 ^ w13518;
	assign w13579 = w13541 ^ w13533;
	assign w13495 = w13527 ^ w43937;
	assign w13538 = w47495 ^ w13495;
	assign w43938 = w13583 ^ w13586;
	assign w13536 = w13584 ^ w43938;
	assign w13492 = w13587 ^ w13536;
	assign w13574 = w47499 ^ w13492;
	assign w13496 = w13522 ^ w43938;
	assign w13580 = w13496 ^ w13521;
	assign w44424 = w25241 ^ w25244;
	assign w25154 = w25180 ^ w44424;
	assign w25238 = w25154 ^ w25179;
	assign w25235 = w25236 ^ w25238;
	assign w25194 = w25242 ^ w44424;
	assign w25150 = w25245 ^ w25194;
	assign w25232 = w47491 ^ w25150;
	assign w44427 = w25241 ^ w25247;
	assign w25153 = w25185 ^ w44427;
	assign w25196 = w47487 ^ w25153;
	assign w25231 = w25236 ^ w25196;
	assign w25230 = w25231 & w25232;
	assign w25228 = w25236 ^ w25230;
	assign w25149 = w25230 ^ w25194;
	assign w25148 = w25230 ^ w25247;
	assign w25143 = w25148 ^ w25244;
	assign w25227 = w25238 & w25228;
	assign w25225 = w25227 ^ w25235;
	assign w44426 = w25227 ^ w25245;
	assign w25219 = w44426 ^ w25197;
	assign w25208 = w25219 & w25260;
	assign w25217 = w25219 & w25256;
	assign w25186 = w47491 ^ w44426;
	assign w25226 = w25186 ^ w25149;
	assign w25216 = w25226 & w25255;
	assign w25207 = w25226 & w25257;
	assign w25229 = w25230 ^ w25238;
	assign w25215 = w25229 & w47492;
	assign w25206 = w25229 & w25261;
	assign w25191 = w44427 ^ w25176;
	assign w25237 = w25199 ^ w25191;
	assign w25234 = w25237 & w25235;
	assign w25233 = w25234 ^ w25196;
	assign w25145 = w25234 ^ w25246;
	assign w25141 = w25145 ^ w25181;
	assign w25144 = w47485 ^ w25141;
	assign w25221 = w25143 ^ w25144;
	assign w25142 = w25234 ^ w25190;
	assign w25140 = w47487 ^ w25141;
	assign w25224 = w25233 & w25225;
	assign w25189 = w25224 ^ w25199;
	assign w25223 = w25189 ^ w25191;
	assign w25147 = w25224 ^ w25248;
	assign w25139 = w25186 ^ w25147;
	assign w25146 = w25176 ^ w25139;
	assign w25222 = w25143 ^ w25146;
	assign w25220 = w25189 ^ w25142;
	assign w25218 = w25139 ^ w25140;
	assign w25214 = w25220 & w25250;
	assign w25213 = w25223 & w25262;
	assign w25212 = w25233 & w25252;
	assign w25156 = w25212 ^ w25213;
	assign w25211 = w25221 & w25253;
	assign w25210 = w25218 & w25251;
	assign w25171 = w25210 ^ w25213;
	assign w25168 = ~w25171;
	assign w25167 = w25210 ^ w25211;
	assign w25209 = w25222 & w25254;
	assign w25205 = w25220 & w25265;
	assign w25187 = w25205 ^ w25209;
	assign w25172 = w25214 ^ w25205;
	assign w25165 = ~w25187;
	assign w25204 = w25223 & w25258;
	assign w25174 = w25212 ^ w25204;
	assign w25203 = w25233 & w25259;
	assign w25164 = w25165 ^ w25203;
	assign w25202 = w25221 & w25264;
	assign w25201 = w25218 & w25266;
	assign w25200 = w25222 & w25263;
	assign w25166 = w25211 ^ w25200;
	assign w25162 = ~w25166;
	assign w44425 = w25201 ^ w25202;
	assign w25183 = w25207 ^ w44425;
	assign w25184 = w25208 ^ w25183;
	assign w25188 = w25216 ^ w25184;
	assign w25157 = w25215 ^ w25188;
	assign w49070 = w25156 ^ w25157;
	assign w7263 = w49070 ^ w7251;
	assign w7517 = w49070 ^ w49074;
	assign w7389 = w7380 ^ w7517;
	assign w48955 = w7389 ^ w7390;
	assign w7359 = w7362 ^ w7517;
	assign w48947 = w7579 ^ w7517;
	assign w47345 = w48947 ^ w1535;
	assign w47337 = w48955 ^ w1543;
	assign w25193 = w25217 ^ w25188;
	assign w25268 = w25193 ^ w25167;
	assign w25170 = w25174 ^ w44425;
	assign w25169 = w25165 ^ w25170;
	assign w25269 = w25168 ^ w25169;
	assign w44428 = w25213 ^ w25214;
	assign w49071 = w44428 ^ w25193;
	assign w7361 = ~w49071;
	assign w7376 = w7361 ^ w49067;
	assign w48965 = w7375 ^ w7376;
	assign w47327 = w48965 ^ w1553;
	assign w7512 = w49071 ^ w49075;
	assign w48948 = w7578 ^ w7512;
	assign w47344 = w48948 ^ w1536;
	assign w7358 = w7516 ^ w7512;
	assign w7386 = w7388 ^ w7512;
	assign w48956 = w7386 ^ w7387;
	assign w47336 = w48956 ^ w1544;
	assign w25195 = w25210 ^ w44428;
	assign w25161 = w25206 ^ w25195;
	assign w25158 = ~w25161;
	assign w25155 = w25211 ^ w25195;
	assign w49072 = w25184 ^ w25155;
	assign w7491 = w49072 ^ w49076;
	assign w7360 = w7491 ^ w7361;
	assign w48972 = w7359 ^ w7360;
	assign w7367 = w7491 ^ w49070;
	assign w47320 = w48972 ^ w1560;
	assign w7382 = w7491 ^ w45262;
	assign w7371 = w7532 ^ w7491;
	assign w48959 = w7382 ^ w7383;
	assign w47333 = w48959 ^ w1547;
	assign w7400 = w7510 ^ w7491;
	assign w48951 = w49068 ^ w7400;
	assign w47341 = w48951 ^ w1539;
	assign w28212 = w47344 ^ w47341;
	assign w13204 = w47336 ^ w47333;
	assign w44429 = w25215 ^ w25217;
	assign w25173 = w44429 ^ w25170;
	assign w25270 = w25172 ^ w25173;
	assign w25160 = w25164 ^ w44429;
	assign w25163 = w25202 ^ w25160;
	assign w25267 = w25162 ^ w25163;
	assign w25159 = w25183 ^ w25160;
	assign w49069 = w25158 ^ w25159;
	assign w7261 = w49069 ^ w49065;
	assign w7522 = w49069 ^ w49073;
	assign w7391 = w7531 ^ w7522;
	assign w7405 = w7522 ^ w45727;
	assign w48954 = w49060 ^ w7391;
	assign w47338 = w48954 ^ w1542;
	assign w13092 = w47337 ^ w47338;
	assign w7366 = w7524 ^ w7522;
	assign w48971 = w7366 ^ w7367;
	assign w47321 = w48971 ^ w1559;
	assign w13581 = w13587 ^ w13539;
	assign w13578 = w13582 & w13581;
	assign w13577 = w13578 ^ w13580;
	assign w13573 = w13578 ^ w13538;
	assign w13576 = w13579 & w13577;
	assign w13487 = w13576 ^ w13588;
	assign w13575 = w13576 ^ w13538;
	assign w13554 = w13575 & w13594;
	assign w13572 = w13573 & w13574;
	assign w13491 = w13572 ^ w13536;
	assign w13490 = w13572 ^ w13589;
	assign w13570 = w13578 ^ w13572;
	assign w13569 = w13580 & w13570;
	assign w13567 = w13569 ^ w13577;
	assign w13566 = w13575 & w13567;
	assign w13489 = w13566 ^ w13590;
	assign w13531 = w13566 ^ w13541;
	assign w13545 = w13575 & w13601;
	assign w13571 = w13572 ^ w13580;
	assign w13557 = w13571 & w47500;
	assign w13548 = w13571 & w13603;
	assign w43941 = w13569 ^ w13587;
	assign w13528 = w47499 ^ w43941;
	assign w13568 = w13528 ^ w13491;
	assign w13558 = w13568 & w13597;
	assign w13481 = w13528 ^ w13489;
	assign w13488 = w13518 ^ w13481;
	assign w13549 = w13568 & w13599;
	assign w13561 = w43941 ^ w13539;
	assign w13559 = w13561 & w13598;
	assign w13550 = w13561 & w13602;
	assign w43940 = w13557 ^ w13559;
	assign w13565 = w13531 ^ w13533;
	assign w13555 = w13565 & w13604;
	assign w13498 = w13554 ^ w13555;
	assign w13546 = w13565 & w13600;
	assign w13516 = w13554 ^ w13546;
	assign w13485 = w13490 ^ w13586;
	assign w13564 = w13485 ^ w13488;
	assign w13551 = w13564 & w13596;
	assign w13483 = w13487 ^ w13523;
	assign w13486 = w47493 ^ w13483;
	assign w13563 = w13485 ^ w13486;
	assign w13482 = w47495 ^ w13483;
	assign w13560 = w13481 ^ w13482;
	assign w13553 = w13563 & w13595;
	assign w13552 = w13560 & w13593;
	assign w13513 = w13552 ^ w13555;
	assign w13510 = ~w13513;
	assign w13509 = w13552 ^ w13553;
	assign w13484 = w13576 ^ w13532;
	assign w13562 = w13531 ^ w13484;
	assign w13556 = w13562 & w13592;
	assign w13547 = w13562 & w13607;
	assign w13529 = w13547 ^ w13551;
	assign w13507 = ~w13529;
	assign w13506 = w13507 ^ w13545;
	assign w13502 = w13506 ^ w43940;
	assign w13514 = w13556 ^ w13547;
	assign w43939 = w13555 ^ w13556;
	assign w13537 = w13552 ^ w43939;
	assign w13497 = w13553 ^ w13537;
	assign w13503 = w13548 ^ w13537;
	assign w13500 = ~w13503;
	assign w13544 = w13563 & w13606;
	assign w13505 = w13544 ^ w13502;
	assign w13543 = w13560 & w13608;
	assign w43534 = w13543 ^ w13544;
	assign w13512 = w13516 ^ w43534;
	assign w13511 = w13507 ^ w13512;
	assign w13611 = w13510 ^ w13511;
	assign w7323 = w45434 ^ w13611;
	assign w49081 = ~w13611;
	assign w7266 = w13611 ^ w45427;
	assign w7572 = w7265 ^ w7266;
	assign w48977 = w7572 ^ w7544;
	assign w47315 = w48977 ^ w1501;
	assign w13515 = w43940 ^ w13512;
	assign w13612 = w13514 ^ w13515;
	assign w13525 = w13549 ^ w43534;
	assign w13526 = w13550 ^ w13525;
	assign w13501 = w13525 ^ w13502;
	assign w49087 = w13526 ^ w13497;
	assign w7341 = w49087 ^ w45433;
	assign w48983 = w7340 ^ w7341;
	assign w13530 = w13558 ^ w13526;
	assign w13535 = w13559 ^ w13530;
	assign w13610 = w13535 ^ w13509;
	assign w49084 = w43939 ^ w13535;
	assign w7321 = w49090 ^ w49084;
	assign w49086 = ~w13610;
	assign w47309 = w48983 ^ w1507;
	assign w18967 = w47309 ^ w47315;
	assign w7497 = w49087 ^ w49091;
	assign w7278 = ~w7497;
	assign w7279 = w7278 ^ w49094;
	assign w7275 = w7278 ^ w49093;
	assign w7493 = w49080 ^ w49087;
	assign w7339 = w7552 ^ w7493;
	assign w7272 = w49084 ^ w49078;
	assign w7570 = w7271 ^ w7272;
	assign w48980 = w7570 ^ w7521;
	assign w47312 = w48980 ^ w1504;
	assign w18966 = w47312 ^ w47309;
	assign w7533 = w49079 ^ w49084;
	assign w7519 = w45433 ^ w49086;
	assign w7319 = w7519 ^ w45643;
	assign w7317 = ~w7319;
	assign w7305 = ~w7533;
	assign w7303 = w7305 ^ w7530;
	assign w7316 = w45441 ^ w13610;
	assign w7330 = w7533 ^ w7515;
	assign w48989 = w45432 ^ w7330;
	assign w47303 = w48989 ^ w1513;
	assign w7301 = w7519 ^ w7515;
	assign w49006 = w45441 ^ w7301;
	assign w47286 = w49006 ^ w1530;
	assign w7328 = w7519 ^ w7490;
	assign w48991 = w49080 ^ w7328;
	assign w47301 = w48991 ^ w1515;
	assign w7300 = w7504 ^ w7493;
	assign w49007 = w49091 ^ w7300;
	assign w47285 = w49007 ^ w1531;
	assign w7344 = w13610 ^ w45432;
	assign w7273 = w7497 ^ w45644;
	assign w7342 = w7343 ^ w7344;
	assign w48982 = ~w7342;
	assign w47310 = w48982 ^ w1506;
	assign w18880 = w47312 ^ w47310;
	assign w49082 = w13500 ^ w13501;
	assign w7548 = w49077 ^ w49082;
	assign w7324 = ~w7548;
	assign w7333 = w7324 ^ w7530;
	assign w7309 = w7548 ^ w7544;
	assign w49002 = w49088 ^ w7309;
	assign w47290 = w49002 ^ w1526;
	assign w31159 = w47285 ^ w47290;
	assign w7322 = w7324 ^ w49092;
	assign w48994 = w7322 ^ w7323;
	assign w47298 = w48994 ^ w1518;
	assign w7277 = ~w49082;
	assign w7352 = w7277 ^ w45426;
	assign w7276 = w49088 ^ w7277;
	assign w48978 = w7351 ^ w7352;
	assign w47314 = w48978 ^ w1502;
	assign w18894 = w47315 ^ w47314;
	assign w18962 = w18966 ^ w18894;
	assign w18968 = w47314 ^ w47312;
	assign w18965 = w47309 ^ w47314;
	assign w7568 = w7275 ^ w7276;
	assign w13499 = w13557 ^ w13530;
	assign w49083 = w13498 ^ w13499;
	assign w7270 = ~w49083;
	assign w7280 = w49089 ^ w7270;
	assign w7567 = w7279 ^ w7280;
	assign w48996 = w7567 ^ w7533;
	assign w47296 = w48996 ^ w1520;
	assign w28080 = w47298 ^ w47296;
	assign w7269 = w7270 ^ w49077;
	assign w7571 = w7268 ^ w7269;
	assign w48979 = w7571 ^ w7530;
	assign w47313 = w48979 ^ w1503;
	assign w18877 = w47315 ^ w47313;
	assign w18879 = w47314 ^ w18877;
	assign w18955 = w47310 ^ w18879;
	assign w18958 = w18877 ^ w18966;
	assign w18854 = w47313 ^ w47314;
	assign w18951 = w18958 & w18962;
	assign w18883 = w18951 ^ w18880;
	assign w18945 = w18966 & w18955;
	assign w18881 = w18945 ^ w18879;
	assign w18887 = w18883 ^ w18881;
	assign w18892 = w47309 ^ w18887;
	assign w7541 = w49078 ^ w49083;
	assign w7308 = ~w7541;
	assign w48995 = w7568 ^ w7541;
	assign w47297 = w48995 ^ w1519;
	assign w27966 = w47297 ^ w47298;
	assign w7331 = w7308 ^ w7521;
	assign w7306 = w7308 ^ w7540;
	assign w13542 = w13564 & w13605;
	assign w13508 = w13553 ^ w13542;
	assign w13504 = ~w13508;
	assign w13609 = w13504 ^ w13505;
	assign w49085 = ~w13609;
	assign w7349 = w13609 ^ w49079;
	assign w7526 = w45432 ^ w49085;
	assign w7320 = w7526 ^ w45642;
	assign w48997 = w7320 ^ w7321;
	assign w47295 = w48997 ^ w1521;
	assign w7318 = w45440 ^ w13609;
	assign w48998 = w7317 ^ w7318;
	assign w47294 = w48998 ^ w1522;
	assign w27992 = w47296 ^ w47294;
	assign w27951 = w27992 ^ w47295;
	assign w7329 = w7526 ^ w7504;
	assign w7302 = w7526 ^ w7521;
	assign w48990 = w45433 ^ w7329;
	assign w47302 = w48990 ^ w1514;
	assign w49005 = w45440 ^ w7302;
	assign w47287 = w49005 ^ w1529;
	assign w31072 = w47287 ^ w47285;
	assign w48981 = w7348 ^ w7349;
	assign w47311 = w48981 ^ w1505;
	assign w18952 = w47311 ^ w18879;
	assign w18878 = w47311 ^ w47309;
	assign w18953 = w18878 ^ w18968;
	assign w18840 = w18880 ^ w18878;
	assign w18956 = w18877 ^ w18840;
	assign w18839 = w18880 ^ w47311;
	assign w18948 = w18967 & w18952;
	assign w18882 = w18948 ^ w18878;
	assign w18944 = w18968 & w18953;
	assign w18853 = w18944 ^ w18945;
	assign w18900 = w18853 ^ w18854;
	assign w18899 = w18900 ^ w18882;
	assign w18943 = w18965 & w18956;
	assign w13206 = w47338 ^ w47336;
	assign w7499 = w49068 ^ w49072;
	assign w7264 = ~w7499;
	assign w7258 = w7499 ^ w45727;
	assign w7262 = w7264 ^ w49075;
	assign w7573 = w7262 ^ w7263;
	assign w48964 = w7573 ^ w7520;
	assign w47328 = w48964 ^ w1552;
	assign w7260 = w7499 ^ w49074;
	assign w7574 = w7260 ^ w7261;
	assign w48963 = w7574 ^ w7524;
	assign w47329 = w48963 ^ w1551;
	assign w7381 = w7532 ^ w7499;
	assign w48960 = w45728 ^ w7381;
	assign w47332 = w48960 ^ w1548;
	assign w7555 = w45426 ^ w49081;
	assign w7313 = w7555 ^ w7552;
	assign w7311 = ~w7313;
	assign w7335 = w7555 ^ w7540;
	assign w48986 = w49077 ^ w7335;
	assign w47306 = w48986 ^ w1510;
	assign w13069 = w47301 ^ w47306;
	assign w48984 = w45427 ^ w7339;
	assign w47308 = w48984 ^ w1508;
	assign w48946 = w7405 ^ w7406;
	assign w47346 = w48946 ^ w1534;
	assign w28214 = w47346 ^ w47344;
	assign w28100 = w47345 ^ w47346;
	assign w28211 = w47341 ^ w47346;
	assign w13203 = w47333 ^ w47338;
	assign w45266 = ~w13612;
	assign w7274 = w45435 ^ w45266;
	assign w7569 = w7273 ^ w7274;
	assign w48993 = w7569 ^ w7555;
	assign w47299 = w48993 ^ w1517;
	assign w27989 = w47299 ^ w47297;
	assign w27991 = w47298 ^ w27989;
	assign w28067 = w47294 ^ w27991;
	assign w28064 = w47295 ^ w27991;
	assign w28006 = w47299 ^ w47298;
	assign w48976 = w45266 ^ w7354;
	assign w47316 = w48976 ^ w1500;
	assign w18957 = w47316 ^ w18958;
	assign w18884 = w47316 ^ w47310;
	assign w18954 = w18884 ^ w18879;
	assign w18961 = w18878 ^ w18884;
	assign w18959 = w18894 ^ w18961;
	assign w18964 = w47311 ^ w18884;
	assign w18960 = w47315 ^ w18964;
	assign w18963 = w47316 ^ w18839;
	assign w18950 = w18959 & w18957;
	assign w18901 = w18944 ^ w18950;
	assign w18942 = w18901 ^ w18892;
	assign w18949 = w47316 & w18963;
	assign w18947 = w18964 & w18960;
	assign w18941 = w18947 ^ w18899;
	assign w18946 = w18961 & w18954;
	assign w18938 = w18942 & w18941;
	assign w7556 = w45427 ^ w45266;
	assign w7325 = w7556 ^ w7497;
	assign w48992 = w45645 ^ w7325;
	assign w47300 = w48992 ^ w1516;
	assign w27996 = w47300 ^ w47294;
	assign w28066 = w27996 ^ w27991;
	assign w28076 = w47295 ^ w27996;
	assign w28072 = w47299 ^ w28076;
	assign w28075 = w47300 ^ w27951;
	assign w28061 = w47300 & w28075;
	assign w28059 = w28076 & w28072;
	assign w7314 = w7556 ^ w7490;
	assign w49000 = w45435 ^ w7314;
	assign w47292 = w49000 ^ w1524;
	assign w31078 = w47292 ^ w47286;
	assign w31155 = w31072 ^ w31078;
	assign w31158 = w47287 ^ w31078;
	assign w7337 = w7556 ^ w7544;
	assign w44160 = w18943 ^ w18946;
	assign w18856 = w18882 ^ w44160;
	assign w18940 = w18856 ^ w18881;
	assign w18937 = w18938 ^ w18940;
	assign w18896 = w18944 ^ w44160;
	assign w18852 = w18947 ^ w18896;
	assign w18934 = w47315 ^ w18852;
	assign w44163 = w18943 ^ w18949;
	assign w18855 = w18887 ^ w44163;
	assign w18898 = w47311 ^ w18855;
	assign w18933 = w18938 ^ w18898;
	assign w18932 = w18933 & w18934;
	assign w18930 = w18938 ^ w18932;
	assign w18851 = w18932 ^ w18896;
	assign w18850 = w18932 ^ w18949;
	assign w18845 = w18850 ^ w18946;
	assign w18929 = w18940 & w18930;
	assign w18927 = w18929 ^ w18937;
	assign w44162 = w18929 ^ w18947;
	assign w18921 = w44162 ^ w18899;
	assign w18910 = w18921 & w18962;
	assign w18919 = w18921 & w18958;
	assign w18888 = w47315 ^ w44162;
	assign w18928 = w18888 ^ w18851;
	assign w18918 = w18928 & w18957;
	assign w18909 = w18928 & w18959;
	assign w18931 = w18932 ^ w18940;
	assign w18917 = w18931 & w47316;
	assign w18908 = w18931 & w18963;
	assign w18893 = w44163 ^ w18878;
	assign w18939 = w18901 ^ w18893;
	assign w18936 = w18939 & w18937;
	assign w18935 = w18936 ^ w18898;
	assign w18847 = w18936 ^ w18948;
	assign w18843 = w18847 ^ w18883;
	assign w18846 = w47309 ^ w18843;
	assign w18923 = w18845 ^ w18846;
	assign w18844 = w18936 ^ w18892;
	assign w18842 = w47311 ^ w18843;
	assign w18926 = w18935 & w18927;
	assign w18891 = w18926 ^ w18901;
	assign w18925 = w18891 ^ w18893;
	assign w18849 = w18926 ^ w18950;
	assign w18841 = w18888 ^ w18849;
	assign w18848 = w18878 ^ w18841;
	assign w18924 = w18845 ^ w18848;
	assign w18922 = w18891 ^ w18844;
	assign w18920 = w18841 ^ w18842;
	assign w18916 = w18922 & w18952;
	assign w18915 = w18925 & w18964;
	assign w18914 = w18935 & w18954;
	assign w18858 = w18914 ^ w18915;
	assign w18913 = w18923 & w18955;
	assign w18912 = w18920 & w18953;
	assign w18873 = w18912 ^ w18915;
	assign w18870 = ~w18873;
	assign w18869 = w18912 ^ w18913;
	assign w18911 = w18924 & w18956;
	assign w18907 = w18922 & w18967;
	assign w18889 = w18907 ^ w18911;
	assign w18874 = w18916 ^ w18907;
	assign w18867 = ~w18889;
	assign w18906 = w18925 & w18960;
	assign w18876 = w18914 ^ w18906;
	assign w18905 = w18935 & w18961;
	assign w18866 = w18867 ^ w18905;
	assign w18904 = w18923 & w18966;
	assign w18903 = w18920 & w18968;
	assign w18902 = w18924 & w18965;
	assign w18868 = w18913 ^ w18902;
	assign w18864 = ~w18868;
	assign w44161 = w18903 ^ w18904;
	assign w18885 = w18909 ^ w44161;
	assign w18886 = w18910 ^ w18885;
	assign w18890 = w18918 ^ w18886;
	assign w18859 = w18917 ^ w18890;
	assign w49262 = w18858 ^ w18859;
	assign w18895 = w18919 ^ w18890;
	assign w18970 = w18895 ^ w18869;
	assign w18872 = w18876 ^ w44161;
	assign w18871 = w18867 ^ w18872;
	assign w18971 = w18870 ^ w18871;
	assign w44164 = w18915 ^ w18916;
	assign w49263 = w44164 ^ w18895;
	assign w18897 = w18912 ^ w44164;
	assign w18863 = w18908 ^ w18897;
	assign w18860 = ~w18863;
	assign w18857 = w18913 ^ w18897;
	assign w49264 = w18886 ^ w18857;
	assign w44165 = w18917 ^ w18919;
	assign w18875 = w44165 ^ w18872;
	assign w18972 = w18874 ^ w18875;
	assign w18862 = w18866 ^ w44165;
	assign w18865 = w18904 ^ w18862;
	assign w18969 = w18864 ^ w18865;
	assign w18861 = w18885 ^ w18862;
	assign w49261 = w18860 ^ w18861;
	assign w45410 = ~w18972;
	assign w45415 = ~w18969;
	assign w45416 = ~w18970;
	assign w7862 = w49264 ^ w45416;
	assign w45417 = ~w18971;
	assign w12982 = w47303 ^ w47301;
	assign w45550 = ~w25268;
	assign w48958 = w45550 ^ w7384;
	assign w7509 = w45262 ^ w45550;
	assign w7372 = w7509 ^ w7492;
	assign w7401 = w7509 ^ w45726;
	assign w48950 = w7401 ^ w7402;
	assign w47342 = w48950 ^ w1538;
	assign w28126 = w47344 ^ w47342;
	assign w48967 = w49076 ^ w7372;
	assign w47325 = w48967 ^ w1555;
	assign w19012 = w47327 ^ w47325;
	assign w19100 = w47328 ^ w47325;
	assign w7356 = w49072 ^ w45550;
	assign w48975 = w7355 ^ w7356;
	assign w47317 = w48975 ^ w1563;
	assign w24996 = w47320 ^ w47317;
	assign w47334 = w48958 ^ w1546;
	assign w13118 = w47336 ^ w47334;
	assign w45551 = ~w25269;
	assign w7379 = w45551 ^ w13343;
	assign w48962 = w7378 ^ w7379;
	assign w47330 = w48962 ^ w1550;
	assign w19102 = w47330 ^ w47328;
	assign w19087 = w19012 ^ w19102;
	assign w18988 = w47329 ^ w47330;
	assign w19099 = w47325 ^ w47330;
	assign w19078 = w19102 & w19087;
	assign w7525 = w45551 ^ w45727;
	assign w7393 = w7532 ^ w7525;
	assign w7368 = w7527 ^ w7525;
	assign w48970 = w49069 ^ w7368;
	assign w47322 = w48970 ^ w1558;
	assign w24998 = w47322 ^ w47320;
	assign w24884 = w47321 ^ w47322;
	assign w24995 = w47317 ^ w47322;
	assign w7392 = w7393 ^ w7394;
	assign w48953 = ~w7392;
	assign w47339 = w48953 ^ w1541;
	assign w13205 = w47333 ^ w47339;
	assign w13115 = w47339 ^ w47337;
	assign w13117 = w47338 ^ w13115;
	assign w13193 = w47334 ^ w13117;
	assign w13183 = w13204 & w13193;
	assign w13119 = w13183 ^ w13117;
	assign w13196 = w13115 ^ w13204;
	assign w7370 = w7491 ^ w45551;
	assign w13132 = w47339 ^ w47338;
	assign w13200 = w13204 ^ w13132;
	assign w13189 = w13196 & w13200;
	assign w13121 = w13189 ^ w13118;
	assign w13125 = w13121 ^ w13119;
	assign w13130 = w47333 ^ w13125;
	assign w48945 = w7580 ^ w7525;
	assign w47347 = w48945 ^ w1533;
	assign w28123 = w47347 ^ w47345;
	assign w28125 = w47346 ^ w28123;
	assign w28201 = w47342 ^ w28125;
	assign w28204 = w28123 ^ w28212;
	assign w28140 = w47347 ^ w47346;
	assign w28208 = w28212 ^ w28140;
	assign w28213 = w47341 ^ w47347;
	assign w28197 = w28204 & w28208;
	assign w28129 = w28197 ^ w28126;
	assign w28191 = w28212 & w28201;
	assign w28127 = w28191 ^ w28125;
	assign w28133 = w28129 ^ w28127;
	assign w28138 = w47341 ^ w28133;
	assign w45552 = ~w25270;
	assign w7259 = w45552 ^ w45263;
	assign w7575 = w7258 ^ w7259;
	assign w48961 = w7575 ^ w7531;
	assign w47331 = w48961 ^ w1549;
	assign w19011 = w47331 ^ w47329;
	assign w19013 = w47330 ^ w19011;
	assign w19086 = w47327 ^ w19013;
	assign w19092 = w19011 ^ w19100;
	assign w19091 = w47332 ^ w19092;
	assign w19028 = w47331 ^ w47330;
	assign w19096 = w19100 ^ w19028;
	assign w19101 = w47325 ^ w47331;
	assign w19085 = w19092 & w19096;
	assign w19082 = w19101 & w19086;
	assign w19016 = w19082 ^ w19012;
	assign w7529 = w45552 ^ w45728;
	assign w7395 = w7529 ^ w7492;
	assign w48952 = w45548 ^ w7395;
	assign w7407 = w7529 ^ w7501;
	assign w48944 = w45263 ^ w7407;
	assign w47348 = w48944 ^ w1532;
	assign w28203 = w47348 ^ w28204;
	assign w28130 = w47348 ^ w47342;
	assign w28200 = w28130 ^ w28125;
	assign w47340 = w48952 ^ w1540;
	assign w13122 = w47340 ^ w47334;
	assign w13195 = w47340 ^ w13196;
	assign w13192 = w13122 ^ w13117;
	assign w7369 = w7531 ^ w7529;
	assign w48968 = w45552 ^ w7371;
	assign w47324 = w48968 ^ w1556;
	assign w48969 = w7369 ^ w7370;
	assign w47323 = w48969 ^ w1557;
	assign w24907 = w47323 ^ w47321;
	assign w24909 = w47322 ^ w24907;
	assign w24988 = w24907 ^ w24996;
	assign w24987 = w47324 ^ w24988;
	assign w24924 = w47323 ^ w47322;
	assign w24992 = w24996 ^ w24924;
	assign w24997 = w47317 ^ w47323;
	assign w24981 = w24988 & w24992;
	assign w45557 = ~w25267;
	assign w7373 = w7510 ^ w45557;
	assign w7507 = w45557 ^ w45733;
	assign w7385 = w7520 ^ w7507;
	assign w48957 = w45553 ^ w7385;
	assign w48966 = w7373 ^ w7374;
	assign w47326 = w48966 ^ w1554;
	assign w19089 = w47326 ^ w19013;
	assign w19014 = w47328 ^ w47326;
	assign w19017 = w19085 ^ w19014;
	assign w19018 = w47332 ^ w47326;
	assign w19088 = w19018 ^ w19013;
	assign w19095 = w19012 ^ w19018;
	assign w19093 = w19028 ^ w19095;
	assign w19098 = w47327 ^ w19018;
	assign w19094 = w47331 ^ w19098;
	assign w18974 = w19014 ^ w19012;
	assign w19090 = w19011 ^ w18974;
	assign w18973 = w19014 ^ w47327;
	assign w19097 = w47332 ^ w18973;
	assign w19084 = w19093 & w19091;
	assign w19035 = w19078 ^ w19084;
	assign w19083 = w47332 & w19097;
	assign w19081 = w19098 & w19094;
	assign w19080 = w19095 & w19088;
	assign w19079 = w19100 & w19089;
	assign w19015 = w19079 ^ w19013;
	assign w19021 = w19017 ^ w19015;
	assign w19026 = w47325 ^ w19021;
	assign w19076 = w19035 ^ w19026;
	assign w18987 = w19078 ^ w19079;
	assign w19034 = w18987 ^ w18988;
	assign w19033 = w19034 ^ w19016;
	assign w19075 = w19081 ^ w19033;
	assign w19077 = w19099 & w19090;
	assign w19072 = w19076 & w19075;
	assign w7403 = w7507 ^ w49075;
	assign w48949 = w7403 ^ w7404;
	assign w47343 = w48949 ^ w1537;
	assign w28198 = w47343 ^ w28125;
	assign w28124 = w47343 ^ w47341;
	assign w28199 = w28124 ^ w28214;
	assign w28207 = w28124 ^ w28130;
	assign w28205 = w28140 ^ w28207;
	assign w28210 = w47343 ^ w28130;
	assign w28206 = w47347 ^ w28210;
	assign w28086 = w28126 ^ w28124;
	assign w28202 = w28123 ^ w28086;
	assign w28085 = w28126 ^ w47343;
	assign w28209 = w47348 ^ w28085;
	assign w28196 = w28205 & w28203;
	assign w28195 = w47348 & w28209;
	assign w28194 = w28213 & w28198;
	assign w28128 = w28194 ^ w28124;
	assign w28193 = w28210 & w28206;
	assign w28192 = w28207 & w28200;
	assign w28190 = w28214 & w28199;
	assign w28147 = w28190 ^ w28196;
	assign w28188 = w28147 ^ w28138;
	assign w28099 = w28190 ^ w28191;
	assign w28146 = w28099 ^ w28100;
	assign w28145 = w28146 ^ w28128;
	assign w28187 = w28193 ^ w28145;
	assign w28189 = w28211 & w28202;
	assign w28184 = w28188 & w28187;
	assign w47335 = w48957 ^ w1545;
	assign w13077 = w13118 ^ w47335;
	assign w13201 = w47340 ^ w13077;
	assign w13116 = w47335 ^ w47333;
	assign w13078 = w13118 ^ w13116;
	assign w13194 = w13115 ^ w13078;
	assign w13181 = w13203 & w13194;
	assign w13191 = w13116 ^ w13206;
	assign w13182 = w13206 & w13191;
	assign w13202 = w47335 ^ w13122;
	assign w13198 = w47339 ^ w13202;
	assign w13190 = w47335 ^ w13117;
	assign w7357 = w7509 ^ w7507;
	assign w48974 = w45546 ^ w7357;
	assign w47318 = w48974 ^ w1562;
	assign w24985 = w47318 ^ w24909;
	assign w24910 = w47320 ^ w47318;
	assign w24913 = w24981 ^ w24910;
	assign w24914 = w47324 ^ w47318;
	assign w24984 = w24914 ^ w24909;
	assign w24975 = w24996 & w24985;
	assign w24911 = w24975 ^ w24909;
	assign w24917 = w24913 ^ w24911;
	assign w24922 = w47317 ^ w24917;
	assign w13185 = w13202 & w13198;
	assign w13187 = w47340 & w13201;
	assign w48973 = w45557 ^ w7358;
	assign w47319 = w48973 ^ w1561;
	assign w24982 = w47319 ^ w24909;
	assign w24908 = w47319 ^ w47317;
	assign w24983 = w24908 ^ w24998;
	assign w24991 = w24908 ^ w24914;
	assign w24989 = w24924 ^ w24991;
	assign w24994 = w47319 ^ w24914;
	assign w24990 = w47323 ^ w24994;
	assign w24870 = w24910 ^ w24908;
	assign w24986 = w24907 ^ w24870;
	assign w24869 = w24910 ^ w47319;
	assign w24993 = w47324 ^ w24869;
	assign w24980 = w24989 & w24987;
	assign w24979 = w47324 & w24993;
	assign w24978 = w24997 & w24982;
	assign w24912 = w24978 ^ w24908;
	assign w24977 = w24994 & w24990;
	assign w24976 = w24991 & w24984;
	assign w24974 = w24998 & w24983;
	assign w24931 = w24974 ^ w24980;
	assign w24972 = w24931 ^ w24922;
	assign w24883 = w24974 ^ w24975;
	assign w24930 = w24883 ^ w24884;
	assign w24929 = w24930 ^ w24912;
	assign w24971 = w24977 ^ w24929;
	assign w24973 = w24995 & w24986;
	assign w24968 = w24972 & w24971;
	assign w13186 = w13205 & w13190;
	assign w13120 = w13186 ^ w13116;
	assign w13091 = w13182 ^ w13183;
	assign w13138 = w13091 ^ w13092;
	assign w13137 = w13138 ^ w13120;
	assign w13179 = w13185 ^ w13137;
	assign w13199 = w13116 ^ w13122;
	assign w13184 = w13199 & w13192;
	assign w13197 = w13132 ^ w13199;
	assign w13188 = w13197 & w13195;
	assign w13139 = w13182 ^ w13188;
	assign w13180 = w13139 ^ w13130;
	assign w13176 = w13180 & w13179;
	assign w43920 = w13181 ^ w13184;
	assign w13094 = w13120 ^ w43920;
	assign w13178 = w13094 ^ w13119;
	assign w13175 = w13176 ^ w13178;
	assign w13134 = w13182 ^ w43920;
	assign w13090 = w13185 ^ w13134;
	assign w13172 = w47339 ^ w13090;
	assign w43923 = w13181 ^ w13187;
	assign w13093 = w13125 ^ w43923;
	assign w13136 = w47335 ^ w13093;
	assign w13171 = w13176 ^ w13136;
	assign w13170 = w13171 & w13172;
	assign w13089 = w13170 ^ w13134;
	assign w13088 = w13170 ^ w13187;
	assign w13168 = w13176 ^ w13170;
	assign w13169 = w13170 ^ w13178;
	assign w13155 = w13169 & w47340;
	assign w13131 = w43923 ^ w13116;
	assign w13177 = w13139 ^ w13131;
	assign w13174 = w13177 & w13175;
	assign w13085 = w13174 ^ w13186;
	assign w13081 = w13085 ^ w13121;
	assign w13080 = w47335 ^ w13081;
	assign w13173 = w13174 ^ w13136;
	assign w13152 = w13173 & w13192;
	assign w13143 = w13173 & w13199;
	assign w13084 = w47333 ^ w13081;
	assign w13082 = w13174 ^ w13130;
	assign w44166 = w19077 ^ w19083;
	assign w19027 = w44166 ^ w19012;
	assign w19073 = w19035 ^ w19027;
	assign w18989 = w19021 ^ w44166;
	assign w19032 = w47327 ^ w18989;
	assign w19067 = w19072 ^ w19032;
	assign w44167 = w19077 ^ w19080;
	assign w19030 = w19078 ^ w44167;
	assign w18986 = w19081 ^ w19030;
	assign w19068 = w47331 ^ w18986;
	assign w19066 = w19067 & w19068;
	assign w19064 = w19072 ^ w19066;
	assign w18985 = w19066 ^ w19030;
	assign w18984 = w19066 ^ w19083;
	assign w18979 = w18984 ^ w19080;
	assign w18990 = w19016 ^ w44167;
	assign w19074 = w18990 ^ w19015;
	assign w19065 = w19066 ^ w19074;
	assign w19071 = w19072 ^ w19074;
	assign w19070 = w19073 & w19071;
	assign w19069 = w19070 ^ w19032;
	assign w18981 = w19070 ^ w19082;
	assign w18977 = w18981 ^ w19017;
	assign w18980 = w47325 ^ w18977;
	assign w19057 = w18979 ^ w18980;
	assign w18978 = w19070 ^ w19026;
	assign w18976 = w47327 ^ w18977;
	assign w19063 = w19074 & w19064;
	assign w19061 = w19063 ^ w19071;
	assign w19060 = w19069 & w19061;
	assign w19025 = w19060 ^ w19035;
	assign w19059 = w19025 ^ w19027;
	assign w18983 = w19060 ^ w19084;
	assign w19056 = w19025 ^ w18978;
	assign w19051 = w19065 & w47332;
	assign w19050 = w19056 & w19086;
	assign w19049 = w19059 & w19098;
	assign w19048 = w19069 & w19088;
	assign w18992 = w19048 ^ w19049;
	assign w19047 = w19057 & w19089;
	assign w19042 = w19065 & w19097;
	assign w19041 = w19056 & w19101;
	assign w19008 = w19050 ^ w19041;
	assign w19040 = w19059 & w19094;
	assign w19010 = w19048 ^ w19040;
	assign w19039 = w19069 & w19095;
	assign w19038 = w19057 & w19100;
	assign w44168 = w19049 ^ w19050;
	assign w44170 = w19063 ^ w19081;
	assign w19022 = w47331 ^ w44170;
	assign w18975 = w19022 ^ w18983;
	assign w18982 = w19012 ^ w18975;
	assign w19058 = w18979 ^ w18982;
	assign w19054 = w18975 ^ w18976;
	assign w19046 = w19054 & w19087;
	assign w19031 = w19046 ^ w44168;
	assign w19007 = w19046 ^ w19049;
	assign w19004 = ~w19007;
	assign w19003 = w19046 ^ w19047;
	assign w18991 = w19047 ^ w19031;
	assign w19045 = w19058 & w19090;
	assign w18997 = w19042 ^ w19031;
	assign w18994 = ~w18997;
	assign w19023 = w19041 ^ w19045;
	assign w19001 = ~w19023;
	assign w19000 = w19001 ^ w19039;
	assign w19037 = w19054 & w19102;
	assign w19036 = w19058 & w19099;
	assign w19002 = w19047 ^ w19036;
	assign w18998 = ~w19002;
	assign w43551 = w19037 ^ w19038;
	assign w19006 = w19010 ^ w43551;
	assign w19005 = w19001 ^ w19006;
	assign w19105 = w19004 ^ w19005;
	assign w19062 = w19022 ^ w18985;
	assign w19052 = w19062 & w19091;
	assign w19043 = w19062 & w19093;
	assign w19019 = w19043 ^ w43551;
	assign w19055 = w44170 ^ w19033;
	assign w19053 = w19055 & w19092;
	assign w19044 = w19055 & w19096;
	assign w19020 = w19044 ^ w19019;
	assign w19024 = w19052 ^ w19020;
	assign w19029 = w19053 ^ w19024;
	assign w49291 = w44168 ^ w19029;
	assign w19104 = w19029 ^ w19003;
	assign w18993 = w19051 ^ w19024;
	assign w49290 = w18992 ^ w18993;
	assign w49292 = w19020 ^ w18991;
	assign w44169 = w19051 ^ w19053;
	assign w19009 = w44169 ^ w19006;
	assign w19106 = w19008 ^ w19009;
	assign w18996 = w19000 ^ w44169;
	assign w18999 = w19038 ^ w18996;
	assign w19103 = w18998 ^ w18999;
	assign w18995 = w19019 ^ w18996;
	assign w49289 = w18994 ^ w18995;
	assign w13083 = w13088 ^ w13184;
	assign w13161 = w13083 ^ w13084;
	assign w13142 = w13161 & w13204;
	assign w44413 = w24973 ^ w24976;
	assign w24886 = w24912 ^ w44413;
	assign w24970 = w24886 ^ w24911;
	assign w24967 = w24968 ^ w24970;
	assign w24926 = w24974 ^ w44413;
	assign w24882 = w24977 ^ w24926;
	assign w24964 = w47323 ^ w24882;
	assign w44416 = w24973 ^ w24979;
	assign w24885 = w24917 ^ w44416;
	assign w24928 = w47319 ^ w24885;
	assign w24963 = w24968 ^ w24928;
	assign w24962 = w24963 & w24964;
	assign w24961 = w24962 ^ w24970;
	assign w24960 = w24968 ^ w24962;
	assign w24881 = w24962 ^ w24926;
	assign w24880 = w24962 ^ w24979;
	assign w24875 = w24880 ^ w24976;
	assign w24959 = w24970 & w24960;
	assign w24957 = w24959 ^ w24967;
	assign w24947 = w24961 & w47324;
	assign w24938 = w24961 & w24993;
	assign w44415 = w24959 ^ w24977;
	assign w24951 = w44415 ^ w24929;
	assign w24949 = w24951 & w24988;
	assign w24940 = w24951 & w24992;
	assign w24918 = w47323 ^ w44415;
	assign w24958 = w24918 ^ w24881;
	assign w24948 = w24958 & w24987;
	assign w24939 = w24958 & w24989;
	assign w24923 = w44416 ^ w24908;
	assign w24969 = w24931 ^ w24923;
	assign w24966 = w24969 & w24967;
	assign w24965 = w24966 ^ w24928;
	assign w24877 = w24966 ^ w24978;
	assign w24873 = w24877 ^ w24913;
	assign w24876 = w47317 ^ w24873;
	assign w24953 = w24875 ^ w24876;
	assign w24874 = w24966 ^ w24922;
	assign w24872 = w47319 ^ w24873;
	assign w24956 = w24965 & w24957;
	assign w24921 = w24956 ^ w24931;
	assign w24955 = w24921 ^ w24923;
	assign w24879 = w24956 ^ w24980;
	assign w24871 = w24918 ^ w24879;
	assign w24878 = w24908 ^ w24871;
	assign w24954 = w24875 ^ w24878;
	assign w24952 = w24921 ^ w24874;
	assign w24950 = w24871 ^ w24872;
	assign w24946 = w24952 & w24982;
	assign w24945 = w24955 & w24994;
	assign w24944 = w24965 & w24984;
	assign w24888 = w24944 ^ w24945;
	assign w24943 = w24953 & w24985;
	assign w24942 = w24950 & w24983;
	assign w24903 = w24942 ^ w24945;
	assign w24900 = ~w24903;
	assign w24899 = w24942 ^ w24943;
	assign w24941 = w24954 & w24986;
	assign w24937 = w24952 & w24997;
	assign w24919 = w24937 ^ w24941;
	assign w24904 = w24946 ^ w24937;
	assign w24897 = ~w24919;
	assign w24936 = w24955 & w24990;
	assign w24906 = w24944 ^ w24936;
	assign w24935 = w24965 & w24991;
	assign w24896 = w24897 ^ w24935;
	assign w24934 = w24953 & w24996;
	assign w24933 = w24950 & w24998;
	assign w24932 = w24954 & w24995;
	assign w24898 = w24943 ^ w24932;
	assign w24894 = ~w24898;
	assign w44414 = w24933 ^ w24934;
	assign w24915 = w24939 ^ w44414;
	assign w24916 = w24940 ^ w24915;
	assign w24920 = w24948 ^ w24916;
	assign w24925 = w24949 ^ w24920;
	assign w25000 = w24925 ^ w24899;
	assign w24889 = w24947 ^ w24920;
	assign w49275 = w24888 ^ w24889;
	assign w24902 = w24906 ^ w44414;
	assign w24901 = w24897 ^ w24902;
	assign w25001 = w24900 ^ w24901;
	assign w44417 = w24945 ^ w24946;
	assign w49276 = w44417 ^ w24925;
	assign w24927 = w24942 ^ w44417;
	assign w24893 = w24938 ^ w24927;
	assign w24890 = ~w24893;
	assign w24887 = w24943 ^ w24927;
	assign w49277 = w24916 ^ w24887;
	assign w7980 = w49264 ^ w49277;
	assign w7731 = w7980 ^ w49275;
	assign w7727 = ~w7980;
	assign w44418 = w24947 ^ w24949;
	assign w24905 = w44418 ^ w24902;
	assign w25002 = w24904 ^ w24905;
	assign w24892 = w24896 ^ w44418;
	assign w24895 = w24934 ^ w24892;
	assign w24999 = w24894 ^ w24895;
	assign w24891 = w24915 ^ w24892;
	assign w49274 = w24890 ^ w24891;
	assign w7728 = w7727 ^ w49274;
	assign w44545 = w28189 ^ w28195;
	assign w28101 = w28133 ^ w44545;
	assign w28144 = w47343 ^ w28101;
	assign w28179 = w28184 ^ w28144;
	assign w28139 = w44545 ^ w28124;
	assign w28185 = w28147 ^ w28139;
	assign w44546 = w28189 ^ w28192;
	assign w28142 = w28190 ^ w44546;
	assign w28098 = w28193 ^ w28142;
	assign w28180 = w47347 ^ w28098;
	assign w28178 = w28179 & w28180;
	assign w28176 = w28184 ^ w28178;
	assign w28097 = w28178 ^ w28142;
	assign w28096 = w28178 ^ w28195;
	assign w28091 = w28096 ^ w28192;
	assign w28102 = w28128 ^ w44546;
	assign w28186 = w28102 ^ w28127;
	assign w28177 = w28178 ^ w28186;
	assign w28183 = w28184 ^ w28186;
	assign w28182 = w28185 & w28183;
	assign w28181 = w28182 ^ w28144;
	assign w28093 = w28182 ^ w28194;
	assign w28089 = w28093 ^ w28129;
	assign w28092 = w47341 ^ w28089;
	assign w28169 = w28091 ^ w28092;
	assign w28090 = w28182 ^ w28138;
	assign w28088 = w47343 ^ w28089;
	assign w28175 = w28186 & w28176;
	assign w28173 = w28175 ^ w28183;
	assign w28172 = w28181 & w28173;
	assign w28137 = w28172 ^ w28147;
	assign w28171 = w28137 ^ w28139;
	assign w28095 = w28172 ^ w28196;
	assign w28168 = w28137 ^ w28090;
	assign w28163 = w28177 & w47348;
	assign w28162 = w28168 & w28198;
	assign w28161 = w28171 & w28210;
	assign w28160 = w28181 & w28200;
	assign w28104 = w28160 ^ w28161;
	assign w28159 = w28169 & w28201;
	assign w28154 = w28177 & w28209;
	assign w28153 = w28168 & w28213;
	assign w28120 = w28162 ^ w28153;
	assign w28152 = w28171 & w28206;
	assign w28122 = w28160 ^ w28152;
	assign w28151 = w28181 & w28207;
	assign w28150 = w28169 & w28212;
	assign w44548 = w28161 ^ w28162;
	assign w44550 = w28175 ^ w28193;
	assign w28167 = w44550 ^ w28145;
	assign w28165 = w28167 & w28204;
	assign w44549 = w28163 ^ w28165;
	assign w28156 = w28167 & w28208;
	assign w28134 = w47347 ^ w44550;
	assign w28174 = w28134 ^ w28097;
	assign w28087 = w28134 ^ w28095;
	assign w28094 = w28124 ^ w28087;
	assign w28170 = w28091 ^ w28094;
	assign w28166 = w28087 ^ w28088;
	assign w28164 = w28174 & w28203;
	assign w28158 = w28166 & w28199;
	assign w28143 = w28158 ^ w44548;
	assign w28119 = w28158 ^ w28161;
	assign w28116 = ~w28119;
	assign w28115 = w28158 ^ w28159;
	assign w28109 = w28154 ^ w28143;
	assign w28106 = ~w28109;
	assign w28103 = w28159 ^ w28143;
	assign w28157 = w28170 & w28202;
	assign w28135 = w28153 ^ w28157;
	assign w28113 = ~w28135;
	assign w28112 = w28113 ^ w28151;
	assign w28108 = w28112 ^ w44549;
	assign w28111 = w28150 ^ w28108;
	assign w28155 = w28174 & w28205;
	assign w28149 = w28166 & w28214;
	assign w28148 = w28170 & w28211;
	assign w28114 = w28159 ^ w28148;
	assign w28110 = ~w28114;
	assign w28215 = w28110 ^ w28111;
	assign w44547 = w28149 ^ w28150;
	assign w28131 = w28155 ^ w44547;
	assign w28107 = w28131 ^ w28108;
	assign w49241 = w28106 ^ w28107;
	assign w28132 = w28156 ^ w28131;
	assign w49244 = w28132 ^ w28103;
	assign w28136 = w28164 ^ w28132;
	assign w28105 = w28163 ^ w28136;
	assign w49242 = w28104 ^ w28105;
	assign w28141 = w28165 ^ w28136;
	assign w28216 = w28141 ^ w28115;
	assign w49243 = w44548 ^ w28141;
	assign w28118 = w28122 ^ w44547;
	assign w28121 = w44549 ^ w28118;
	assign w28218 = w28120 ^ w28121;
	assign w28117 = w28113 ^ w28118;
	assign w28217 = w28116 ^ w28117;
	assign w13167 = w13178 & w13168;
	assign w13165 = w13167 ^ w13175;
	assign w13164 = w13173 & w13165;
	assign w13129 = w13164 ^ w13139;
	assign w13163 = w13129 ^ w13131;
	assign w13153 = w13163 & w13202;
	assign w13096 = w13152 ^ w13153;
	assign w13160 = w13129 ^ w13082;
	assign w13154 = w13160 & w13190;
	assign w13145 = w13160 & w13205;
	assign w13112 = w13154 ^ w13145;
	assign w13144 = w13163 & w13198;
	assign w13114 = w13152 ^ w13144;
	assign w43922 = w13167 ^ w13185;
	assign w13159 = w43922 ^ w13137;
	assign w13148 = w13159 & w13200;
	assign w13157 = w13159 & w13196;
	assign w13126 = w47339 ^ w43922;
	assign w13166 = w13126 ^ w13089;
	assign w13156 = w13166 & w13195;
	assign w13147 = w13166 & w13197;
	assign w43924 = w13153 ^ w13154;
	assign w43925 = w13155 ^ w13157;
	assign w13087 = w13164 ^ w13188;
	assign w13079 = w13126 ^ w13087;
	assign w13086 = w13116 ^ w13079;
	assign w13162 = w13083 ^ w13086;
	assign w13140 = w13162 & w13203;
	assign w13149 = w13162 & w13194;
	assign w13127 = w13145 ^ w13149;
	assign w13105 = ~w13127;
	assign w13104 = w13105 ^ w13143;
	assign w13100 = w13104 ^ w43925;
	assign w13103 = w13142 ^ w13100;
	assign w13158 = w13079 ^ w13080;
	assign w13150 = w13158 & w13191;
	assign w13135 = w13150 ^ w43924;
	assign w13111 = w13150 ^ w13153;
	assign w13108 = ~w13111;
	assign w13141 = w13158 & w13206;
	assign w43921 = w13141 ^ w13142;
	assign w13123 = w13147 ^ w43921;
	assign w13124 = w13148 ^ w13123;
	assign w13128 = w13156 ^ w13124;
	assign w13097 = w13155 ^ w13128;
	assign w49303 = w13096 ^ w13097;
	assign w13133 = w13157 ^ w13128;
	assign w49304 = w43924 ^ w13133;
	assign w13099 = w13123 ^ w13100;
	assign w13110 = w13114 ^ w43921;
	assign w13113 = w43925 ^ w13110;
	assign w13210 = w13112 ^ w13113;
	assign w13109 = w13105 ^ w13110;
	assign w13209 = w13108 ^ w13109;
	assign w13151 = w13161 & w13193;
	assign w13107 = w13150 ^ w13151;
	assign w13095 = w13151 ^ w13135;
	assign w49305 = w13124 ^ w13095;
	assign w13208 = w13133 ^ w13107;
	assign w13106 = w13151 ^ w13140;
	assign w13102 = ~w13106;
	assign w13207 = w13102 ^ w13103;
	assign w45258 = ~w13209;
	assign w45259 = ~w13210;
	assign w45264 = ~w13207;
	assign w7937 = w45264 ^ w49304;
	assign w45265 = ~w13208;
	assign w45414 = ~w19106;
	assign w45419 = ~w19103;
	assign w45420 = ~w19104;
	assign w45421 = ~w19105;
	assign w45542 = ~w25000;
	assign w7989 = w45416 ^ w45542;
	assign w45543 = ~w25001;
	assign w45544 = ~w25002;
	assign w7725 = w7727 ^ w45544;
	assign w45549 = ~w24999;
	assign w7881 = w45549 ^ w45415;
	assign w45634 = ~w28216;
	assign w45635 = ~w28217;
	assign w7767 = w45635 ^ w45409;
	assign w7948 = w45635 ^ w7770;
	assign w45636 = ~w28218;
	assign w7763 = w18703 ^ w45636;
	assign w45641 = ~w28215;
	assign w13146 = w13169 & w13201;
	assign w13101 = w13146 ^ w13135;
	assign w13098 = ~w13101;
	assign w49302 = w13098 ^ w13099;
	assign w7722 = w49303 ^ w49302;
	assign w12988 = w47308 ^ w47302;
	assign w13065 = w12982 ^ w12988;
	assign w13068 = w47303 ^ w12988;
	assign w45893 = ~w7493;
	assign w7334 = w45893 ^ w49078;
	assign w48987 = w7333 ^ w7334;
	assign w47305 = w48987 ^ w1511;
	assign w12958 = w47305 ^ w47306;
	assign w7332 = w45893 ^ w49079;
	assign w7315 = w45893 ^ w49095;
	assign w48988 = w7331 ^ w7332;
	assign w47304 = w48988 ^ w1512;
	assign w13072 = w47306 ^ w47304;
	assign w13057 = w12982 ^ w13072;
	assign w48999 = w7315 ^ w7316;
	assign w47293 = w48999 ^ w1523;
	assign w27990 = w47295 ^ w47293;
	assign w28065 = w27990 ^ w28080;
	assign w28078 = w47296 ^ w47293;
	assign w28074 = w28078 ^ w28006;
	assign w28073 = w27990 ^ w27996;
	assign w28071 = w28006 ^ w28073;
	assign w28070 = w27989 ^ w28078;
	assign w28069 = w47300 ^ w28070;
	assign w27952 = w27992 ^ w27990;
	assign w28068 = w27989 ^ w27952;
	assign w28079 = w47293 ^ w47299;
	assign w28077 = w47293 ^ w47298;
	assign w28063 = w28070 & w28074;
	assign w27995 = w28063 ^ w27992;
	assign w28062 = w28071 & w28069;
	assign w28060 = w28079 & w28064;
	assign w27994 = w28060 ^ w27990;
	assign w28058 = w28073 & w28066;
	assign w28057 = w28078 & w28067;
	assign w27993 = w28057 ^ w27991;
	assign w27999 = w27995 ^ w27993;
	assign w28004 = w47293 ^ w27999;
	assign w28056 = w28080 & w28065;
	assign w28013 = w28056 ^ w28062;
	assign w28054 = w28013 ^ w28004;
	assign w27965 = w28056 ^ w28057;
	assign w28012 = w27965 ^ w27966;
	assign w28011 = w28012 ^ w27994;
	assign w28053 = w28059 ^ w28011;
	assign w28055 = w28077 & w28068;
	assign w28050 = w28054 & w28053;
	assign w7338 = w45893 ^ w45426;
	assign w7336 = w7337 ^ w7338;
	assign w48985 = ~w7336;
	assign w47307 = w48985 ^ w1509;
	assign w13071 = w47301 ^ w47307;
	assign w13064 = w47307 ^ w13068;
	assign w13051 = w13068 & w13064;
	assign w12998 = w47307 ^ w47306;
	assign w12984 = w47304 ^ w47302;
	assign w12943 = w12984 ^ w47303;
	assign w12944 = w12984 ^ w12982;
	assign w13067 = w47308 ^ w12943;
	assign w13063 = w12998 ^ w13065;
	assign w13070 = w47304 ^ w47301;
	assign w44540 = w28055 ^ w28061;
	assign w28005 = w44540 ^ w27990;
	assign w28051 = w28013 ^ w28005;
	assign w27967 = w27999 ^ w44540;
	assign w28010 = w47295 ^ w27967;
	assign w28045 = w28050 ^ w28010;
	assign w44541 = w28055 ^ w28058;
	assign w28008 = w28056 ^ w44541;
	assign w27964 = w28059 ^ w28008;
	assign w28046 = w47299 ^ w27964;
	assign w28044 = w28045 & w28046;
	assign w27963 = w28044 ^ w28008;
	assign w27962 = w28044 ^ w28061;
	assign w27957 = w27962 ^ w28058;
	assign w28042 = w28050 ^ w28044;
	assign w27968 = w27994 ^ w44541;
	assign w28052 = w27968 ^ w27993;
	assign w28043 = w28044 ^ w28052;
	assign w28049 = w28050 ^ w28052;
	assign w28048 = w28051 & w28049;
	assign w28047 = w28048 ^ w28010;
	assign w27959 = w28048 ^ w28060;
	assign w27955 = w27959 ^ w27995;
	assign w27958 = w47293 ^ w27955;
	assign w28035 = w27957 ^ w27958;
	assign w27956 = w28048 ^ w28004;
	assign w27954 = w47295 ^ w27955;
	assign w28041 = w28052 & w28042;
	assign w28039 = w28041 ^ w28049;
	assign w28038 = w28047 & w28039;
	assign w28003 = w28038 ^ w28013;
	assign w28037 = w28003 ^ w28005;
	assign w27961 = w28038 ^ w28062;
	assign w28034 = w28003 ^ w27956;
	assign w28029 = w28043 & w47300;
	assign w28028 = w28034 & w28064;
	assign w28027 = w28037 & w28076;
	assign w28026 = w28047 & w28066;
	assign w27970 = w28026 ^ w28027;
	assign w28025 = w28035 & w28067;
	assign w28020 = w28043 & w28075;
	assign w28019 = w28034 & w28079;
	assign w27986 = w28028 ^ w28019;
	assign w28018 = w28037 & w28072;
	assign w27988 = w28026 ^ w28018;
	assign w28017 = w28047 & w28073;
	assign w28016 = w28035 & w28078;
	assign w44542 = w28027 ^ w28028;
	assign w44544 = w28041 ^ w28059;
	assign w28000 = w47299 ^ w44544;
	assign w28040 = w28000 ^ w27963;
	assign w28021 = w28040 & w28071;
	assign w28030 = w28040 & w28069;
	assign w27953 = w28000 ^ w27961;
	assign w27960 = w27990 ^ w27953;
	assign w28036 = w27957 ^ w27960;
	assign w28023 = w28036 & w28068;
	assign w28001 = w28019 ^ w28023;
	assign w27979 = ~w28001;
	assign w27978 = w27979 ^ w28017;
	assign w28032 = w27953 ^ w27954;
	assign w28015 = w28032 & w28080;
	assign w28014 = w28036 & w28077;
	assign w27980 = w28025 ^ w28014;
	assign w27976 = ~w27980;
	assign w43579 = w28015 ^ w28016;
	assign w27997 = w28021 ^ w43579;
	assign w27984 = w27988 ^ w43579;
	assign w27983 = w27979 ^ w27984;
	assign w28024 = w28032 & w28065;
	assign w27981 = w28024 ^ w28025;
	assign w28009 = w28024 ^ w44542;
	assign w27975 = w28020 ^ w28009;
	assign w27972 = ~w27975;
	assign w27969 = w28025 ^ w28009;
	assign w27985 = w28024 ^ w28027;
	assign w27982 = ~w27985;
	assign w28083 = w27982 ^ w27983;
	assign w28033 = w44544 ^ w28011;
	assign w28031 = w28033 & w28070;
	assign w28022 = w28033 & w28074;
	assign w27998 = w28022 ^ w27997;
	assign w28002 = w28030 ^ w27998;
	assign w28007 = w28031 ^ w28002;
	assign w49308 = w44542 ^ w28007;
	assign w28082 = w28007 ^ w27981;
	assign w27971 = w28029 ^ w28002;
	assign w49307 = w27970 ^ w27971;
	assign w7775 = w49308 ^ w49307;
	assign w49309 = w27998 ^ w27969;
	assign w7987 = w49303 ^ w49307;
	assign w7982 = w49305 ^ w49309;
	assign w44543 = w28029 ^ w28031;
	assign w27987 = w44543 ^ w27984;
	assign w28084 = w27986 ^ w27987;
	assign w27974 = w27978 ^ w44543;
	assign w27977 = w28016 ^ w27974;
	assign w28081 = w27976 ^ w27977;
	assign w27973 = w27997 ^ w27974;
	assign w49306 = w27972 ^ w27973;
	assign w7721 = w7982 ^ w49306;
	assign w8061 = w7721 ^ w7722;
	assign w13053 = w47308 & w13067;
	assign w13048 = w13072 & w13057;
	assign w12981 = w47307 ^ w47305;
	assign w13060 = w12981 ^ w12944;
	assign w13047 = w13069 & w13060;
	assign w13062 = w12981 ^ w13070;
	assign w13061 = w47308 ^ w13062;
	assign w13054 = w13063 & w13061;
	assign w13005 = w13048 ^ w13054;
	assign w12983 = w47306 ^ w12981;
	assign w13056 = w47303 ^ w12983;
	assign w13058 = w12988 ^ w12983;
	assign w13052 = w13071 & w13056;
	assign w13050 = w13065 & w13058;
	assign w13059 = w47302 ^ w12983;
	assign w13049 = w13070 & w13059;
	assign w12957 = w13048 ^ w13049;
	assign w13004 = w12957 ^ w12958;
	assign w43915 = w13047 ^ w13050;
	assign w13000 = w13048 ^ w43915;
	assign w12956 = w13051 ^ w13000;
	assign w13038 = w47307 ^ w12956;
	assign w12985 = w13049 ^ w12983;
	assign w12986 = w13052 ^ w12982;
	assign w12960 = w12986 ^ w43915;
	assign w13044 = w12960 ^ w12985;
	assign w13003 = w13004 ^ w12986;
	assign w13045 = w13051 ^ w13003;
	assign w45630 = ~w28082;
	assign w7934 = w45630 ^ w45265;
	assign w45631 = ~w28083;
	assign w7941 = w45631 ^ w45258;
	assign w45632 = ~w28084;
	assign w7720 = w45632 ^ w45259;
	assign w45637 = ~w28081;
	assign w7923 = w45630 ^ w45637;
	assign w7992 = w45264 ^ w45637;
	assign w7963 = ~w7992;
	assign w43914 = w13047 ^ w13053;
	assign w12997 = w43914 ^ w12982;
	assign w13043 = w13005 ^ w12997;
	assign w13066 = w13070 ^ w12998;
	assign w13055 = w13062 & w13066;
	assign w12987 = w13055 ^ w12984;
	assign w12991 = w12987 ^ w12985;
	assign w12996 = w47301 ^ w12991;
	assign w12959 = w12991 ^ w43914;
	assign w13002 = w47303 ^ w12959;
	assign w13046 = w13005 ^ w12996;
	assign w13042 = w13046 & w13045;
	assign w13037 = w13042 ^ w13002;
	assign w13036 = w13037 & w13038;
	assign w13041 = w13042 ^ w13044;
	assign w12955 = w13036 ^ w13000;
	assign w12954 = w13036 ^ w13053;
	assign w12949 = w12954 ^ w13050;
	assign w13040 = w13043 & w13041;
	assign w12951 = w13040 ^ w13052;
	assign w12948 = w13040 ^ w12996;
	assign w12947 = w12951 ^ w12987;
	assign w12950 = w47301 ^ w12947;
	assign w13027 = w12949 ^ w12950;
	assign w13017 = w13027 & w13059;
	assign w13008 = w13027 & w13070;
	assign w12946 = w47303 ^ w12947;
	assign w13039 = w13040 ^ w13002;
	assign w13018 = w13039 & w13058;
	assign w13009 = w13039 & w13065;
	assign w13035 = w13036 ^ w13044;
	assign w13021 = w13035 & w47308;
	assign w13012 = w13035 & w13067;
	assign w13034 = w13042 ^ w13036;
	assign w13033 = w13044 & w13034;
	assign w13031 = w13033 ^ w13041;
	assign w13030 = w13039 & w13031;
	assign w12995 = w13030 ^ w13005;
	assign w12953 = w13030 ^ w13054;
	assign w13026 = w12995 ^ w12948;
	assign w13020 = w13026 & w13056;
	assign w13011 = w13026 & w13071;
	assign w12978 = w13020 ^ w13011;
	assign w43919 = w13033 ^ w13051;
	assign w13025 = w43919 ^ w13003;
	assign w13023 = w13025 & w13062;
	assign w43918 = w13021 ^ w13023;
	assign w13014 = w13025 & w13066;
	assign w12992 = w47307 ^ w43919;
	assign w13032 = w12992 ^ w12955;
	assign w13013 = w13032 & w13063;
	assign w13022 = w13032 & w13061;
	assign w12945 = w12992 ^ w12953;
	assign w12952 = w12982 ^ w12945;
	assign w13028 = w12949 ^ w12952;
	assign w13006 = w13028 & w13069;
	assign w13015 = w13028 & w13060;
	assign w12972 = w13017 ^ w13006;
	assign w12968 = ~w12972;
	assign w13024 = w12945 ^ w12946;
	assign w13016 = w13024 & w13057;
	assign w12973 = w13016 ^ w13017;
	assign w13007 = w13024 & w13072;
	assign w12993 = w13011 ^ w13015;
	assign w12971 = ~w12993;
	assign w12970 = w12971 ^ w13009;
	assign w12966 = w12970 ^ w43918;
	assign w12969 = w13008 ^ w12966;
	assign w13073 = w12968 ^ w12969;
	assign w49248 = ~w13073;
	assign w7901 = w45407 ^ w13073;
	assign w8026 = w45641 ^ w49248;
	assign w43916 = w13007 ^ w13008;
	assign w12989 = w13013 ^ w43916;
	assign w12965 = w12989 ^ w12966;
	assign w12990 = w13014 ^ w12989;
	assign w12994 = w13022 ^ w12990;
	assign w12963 = w13021 ^ w12994;
	assign w12999 = w13023 ^ w12994;
	assign w13074 = w12999 ^ w12973;
	assign w7899 = w45408 ^ w13074;
	assign w49249 = ~w13074;
	assign w8024 = w45634 ^ w49249;
	assign w13029 = w12995 ^ w12997;
	assign w13019 = w13029 & w13068;
	assign w12977 = w13016 ^ w13019;
	assign w12974 = ~w12977;
	assign w12962 = w13018 ^ w13019;
	assign w49246 = w12962 ^ w12963;
	assign w7761 = w49253 ^ w49246;
	assign w13010 = w13029 & w13064;
	assign w12980 = w13018 ^ w13010;
	assign w12976 = w12980 ^ w43916;
	assign w12975 = w12971 ^ w12976;
	assign w13075 = w12974 ^ w12975;
	assign w8038 = w49242 ^ w49246;
	assign w12979 = w43918 ^ w12976;
	assign w13076 = w12978 ^ w12979;
	assign w7920 = ~w8038;
	assign w43917 = w13019 ^ w13020;
	assign w13001 = w13016 ^ w43917;
	assign w12967 = w13012 ^ w13001;
	assign w12961 = w13017 ^ w13001;
	assign w49250 = w12990 ^ w12961;
	assign w7975 = w49250 ^ w49255;
	assign w7909 = ~w7975;
	assign w7974 = w49244 ^ w49250;
	assign w7764 = w7974 ^ w49242;
	assign w12964 = ~w12967;
	assign w49245 = w12964 ^ w12965;
	assign w8013 = w49245 ^ w49252;
	assign w7896 = ~w8013;
	assign w7894 = w7896 ^ w49241;
	assign w7765 = w49241 ^ w49245;
	assign w8043 = w7764 ^ w7765;
	assign w7907 = w8038 ^ w7896;
	assign w49247 = w43917 ^ w12999;
	assign w7903 = w49254 ^ w49247;
	assign w8029 = w49243 ^ w49247;
	assign w45260 = ~w13075;
	assign w8015 = w45260 ^ w49251;
	assign w7913 = w7909 ^ w45260;
	assign w45261 = ~w13076;
	assign w8014 = w45261 ^ w45409;
	assign w45916 = ~w7490;
	assign w7304 = w45916 ^ w49090;
	assign w49004 = w7303 ^ w7304;
	assign w47288 = w49004 ^ w1528;
	assign w31074 = w47288 ^ w47286;
	assign w31160 = w47288 ^ w47285;
	assign w31162 = w47290 ^ w47288;
	assign w31147 = w31072 ^ w31162;
	assign w31034 = w31074 ^ w31072;
	assign w31033 = w31074 ^ w47287;
	assign w31157 = w47292 ^ w31033;
	assign w31143 = w47292 & w31157;
	assign w31138 = w31162 & w31147;
	assign w7312 = w45916 ^ w45434;
	assign w49001 = w7311 ^ w7312;
	assign w47291 = w49001 ^ w1525;
	assign w31154 = w47291 ^ w31158;
	assign w31088 = w47291 ^ w47290;
	assign w31153 = w31088 ^ w31155;
	assign w31156 = w31160 ^ w31088;
	assign w31161 = w47285 ^ w47291;
	assign w31141 = w31158 & w31154;
	assign w7307 = w45916 ^ w49089;
	assign w49003 = w7306 ^ w7307;
	assign w47289 = w49003 ^ w1527;
	assign w31071 = w47291 ^ w47289;
	assign w31073 = w47290 ^ w31071;
	assign w31149 = w47286 ^ w31073;
	assign w31146 = w47287 ^ w31073;
	assign w31148 = w31078 ^ w31073;
	assign w31152 = w31071 ^ w31160;
	assign w31151 = w47292 ^ w31152;
	assign w31048 = w47289 ^ w47290;
	assign w31150 = w31071 ^ w31034;
	assign w31145 = w31152 & w31156;
	assign w31077 = w31145 ^ w31074;
	assign w31144 = w31153 & w31151;
	assign w31095 = w31138 ^ w31144;
	assign w31142 = w31161 & w31146;
	assign w31076 = w31142 ^ w31072;
	assign w31140 = w31155 & w31148;
	assign w31139 = w31160 & w31149;
	assign w31075 = w31139 ^ w31073;
	assign w31081 = w31077 ^ w31075;
	assign w31086 = w47285 ^ w31081;
	assign w31136 = w31095 ^ w31086;
	assign w31047 = w31138 ^ w31139;
	assign w31094 = w31047 ^ w31048;
	assign w31093 = w31094 ^ w31076;
	assign w31135 = w31141 ^ w31093;
	assign w31137 = w31159 & w31150;
	assign w31132 = w31136 & w31135;
	assign w44671 = w31137 ^ w31143;
	assign w31049 = w31081 ^ w44671;
	assign w31092 = w47287 ^ w31049;
	assign w31127 = w31132 ^ w31092;
	assign w31087 = w44671 ^ w31072;
	assign w31133 = w31095 ^ w31087;
	assign w44672 = w31137 ^ w31140;
	assign w31090 = w31138 ^ w44672;
	assign w31046 = w31141 ^ w31090;
	assign w31128 = w47291 ^ w31046;
	assign w31126 = w31127 & w31128;
	assign w31045 = w31126 ^ w31090;
	assign w31124 = w31132 ^ w31126;
	assign w31044 = w31126 ^ w31143;
	assign w31039 = w31044 ^ w31140;
	assign w31050 = w31076 ^ w44672;
	assign w31134 = w31050 ^ w31075;
	assign w31125 = w31126 ^ w31134;
	assign w31131 = w31132 ^ w31134;
	assign w31130 = w31133 & w31131;
	assign w31129 = w31130 ^ w31092;
	assign w31041 = w31130 ^ w31142;
	assign w31037 = w31041 ^ w31077;
	assign w31040 = w47285 ^ w31037;
	assign w31117 = w31039 ^ w31040;
	assign w31038 = w31130 ^ w31086;
	assign w31036 = w47287 ^ w31037;
	assign w31123 = w31134 & w31124;
	assign w31121 = w31123 ^ w31131;
	assign w31120 = w31129 & w31121;
	assign w31085 = w31120 ^ w31095;
	assign w31119 = w31085 ^ w31087;
	assign w31043 = w31120 ^ w31144;
	assign w31116 = w31085 ^ w31038;
	assign w31111 = w31125 & w47292;
	assign w31110 = w31116 & w31146;
	assign w31109 = w31119 & w31158;
	assign w31108 = w31129 & w31148;
	assign w31052 = w31108 ^ w31109;
	assign w31107 = w31117 & w31149;
	assign w31102 = w31125 & w31157;
	assign w31101 = w31116 & w31161;
	assign w31068 = w31110 ^ w31101;
	assign w31100 = w31119 & w31154;
	assign w31070 = w31108 ^ w31100;
	assign w31099 = w31129 & w31155;
	assign w31098 = w31117 & w31160;
	assign w44674 = w31109 ^ w31110;
	assign w44676 = w31123 ^ w31141;
	assign w31115 = w44676 ^ w31093;
	assign w31113 = w31115 & w31152;
	assign w44675 = w31111 ^ w31113;
	assign w31104 = w31115 & w31156;
	assign w31082 = w47291 ^ w44676;
	assign w31122 = w31082 ^ w31045;
	assign w31035 = w31082 ^ w31043;
	assign w31042 = w31072 ^ w31035;
	assign w31118 = w31039 ^ w31042;
	assign w31114 = w31035 ^ w31036;
	assign w31112 = w31122 & w31151;
	assign w31106 = w31114 & w31147;
	assign w31091 = w31106 ^ w44674;
	assign w31067 = w31106 ^ w31109;
	assign w31064 = ~w31067;
	assign w31063 = w31106 ^ w31107;
	assign w31057 = w31102 ^ w31091;
	assign w31054 = ~w31057;
	assign w31051 = w31107 ^ w31091;
	assign w31105 = w31118 & w31150;
	assign w31083 = w31101 ^ w31105;
	assign w31061 = ~w31083;
	assign w31060 = w31061 ^ w31099;
	assign w31056 = w31060 ^ w44675;
	assign w31059 = w31098 ^ w31056;
	assign w31103 = w31122 & w31153;
	assign w31097 = w31114 & w31162;
	assign w31096 = w31118 & w31159;
	assign w31062 = w31107 ^ w31096;
	assign w31058 = ~w31062;
	assign w31163 = w31058 ^ w31059;
	assign w44673 = w31097 ^ w31098;
	assign w31079 = w31103 ^ w44673;
	assign w31055 = w31079 ^ w31056;
	assign w49293 = w31054 ^ w31055;
	assign w31080 = w31104 ^ w31079;
	assign w49296 = w31080 ^ w31051;
	assign w31084 = w31112 ^ w31080;
	assign w31053 = w31111 ^ w31084;
	assign w49294 = w31052 ^ w31053;
	assign w31089 = w31113 ^ w31084;
	assign w31164 = w31089 ^ w31063;
	assign w8019 = w49289 ^ w49293;
	assign w7832 = ~w8019;
	assign w7969 = w49292 ^ w49296;
	assign w8009 = w49290 ^ w49294;
	assign w49295 = w44674 ^ w31089;
	assign w8000 = w49291 ^ w49295;
	assign w31066 = w31070 ^ w44673;
	assign w31069 = w44675 ^ w31066;
	assign w31166 = w31068 ^ w31069;
	assign w31065 = w31061 ^ w31066;
	assign w31165 = w31064 ^ w31065;
	assign w45714 = ~w31165;
	assign w7830 = w7832 ^ w45714;
	assign w8023 = w45421 ^ w45714;
	assign w45715 = ~w31166;
	assign w8031 = w45414 ^ w45715;
	assign w45720 = ~w31163;
	assign w7994 = w45419 ^ w45720;
	assign w7829 = w7994 ^ w49295;
	assign w7827 = ~w7829;
	assign w45721 = ~w31164;
	assign w7819 = w7969 ^ w45721;
	assign w7983 = w45420 ^ w45721;
	assign w7822 = w7983 ^ w45720;
	assign w45917 = ~w7489;
	assign w7477 = w45917 ^ w45442;
	assign w7475 = w7476 ^ w7477;
	assign w49017 = ~w7475;
	assign w7472 = w45917 ^ w49106;
	assign w49019 = w7471 ^ w7472;
	assign w47275 = w49017 ^ w1478;
	assign w34102 = w47275 ^ w34106;
	assign w34036 = w47275 ^ w47274;
	assign w34101 = w34036 ^ w34103;
	assign w34109 = w47269 ^ w47275;
	assign w34089 = w34106 & w34102;
	assign w47273 = w49019 ^ w1480;
	assign w34019 = w47275 ^ w47273;
	assign w34021 = w47274 ^ w34019;
	assign w34097 = w47270 ^ w34021;
	assign w34094 = w47271 ^ w34021;
	assign w34096 = w34026 ^ w34021;
	assign w33996 = w47273 ^ w47274;
	assign w34090 = w34109 & w34094;
	assign w34024 = w34090 ^ w34020;
	assign w34088 = w34103 & w34096;
	assign w7292 = w45917 ^ w49097;
	assign w7561 = w7292 ^ w7293;
	assign w49020 = w7561 ^ w7505;
	assign w47272 = w49020 ^ w1481;
	assign w34022 = w47272 ^ w47270;
	assign w34108 = w47272 ^ w47269;
	assign w34104 = w34108 ^ w34036;
	assign w34100 = w34019 ^ w34108;
	assign w34099 = w47276 ^ w34100;
	assign w34110 = w47274 ^ w47272;
	assign w34095 = w34020 ^ w34110;
	assign w33982 = w34022 ^ w34020;
	assign w34098 = w34019 ^ w33982;
	assign w33981 = w34022 ^ w47271;
	assign w34105 = w47276 ^ w33981;
	assign w34093 = w34100 & w34104;
	assign w34025 = w34093 ^ w34022;
	assign w34092 = w34101 & w34099;
	assign w34091 = w47276 & w34105;
	assign w34087 = w34108 & w34097;
	assign w34023 = w34087 ^ w34021;
	assign w34029 = w34025 ^ w34023;
	assign w34034 = w47269 ^ w34029;
	assign w34086 = w34110 & w34095;
	assign w34043 = w34086 ^ w34092;
	assign w34084 = w34043 ^ w34034;
	assign w33995 = w34086 ^ w34087;
	assign w34042 = w33995 ^ w33996;
	assign w34041 = w34042 ^ w34024;
	assign w34083 = w34089 ^ w34041;
	assign w34085 = w34107 & w34098;
	assign w34080 = w34084 & w34083;
	assign w44794 = w34085 ^ w34091;
	assign w33997 = w34029 ^ w44794;
	assign w34040 = w47271 ^ w33997;
	assign w34075 = w34080 ^ w34040;
	assign w34035 = w44794 ^ w34020;
	assign w34081 = w34043 ^ w34035;
	assign w44795 = w34085 ^ w34088;
	assign w34038 = w34086 ^ w44795;
	assign w33994 = w34089 ^ w34038;
	assign w34076 = w47275 ^ w33994;
	assign w34074 = w34075 & w34076;
	assign w33993 = w34074 ^ w34038;
	assign w34072 = w34080 ^ w34074;
	assign w33992 = w34074 ^ w34091;
	assign w33987 = w33992 ^ w34088;
	assign w33998 = w34024 ^ w44795;
	assign w34082 = w33998 ^ w34023;
	assign w34073 = w34074 ^ w34082;
	assign w34079 = w34080 ^ w34082;
	assign w34078 = w34081 & w34079;
	assign w34077 = w34078 ^ w34040;
	assign w33989 = w34078 ^ w34090;
	assign w33985 = w33989 ^ w34025;
	assign w33988 = w47269 ^ w33985;
	assign w34065 = w33987 ^ w33988;
	assign w33986 = w34078 ^ w34034;
	assign w33984 = w47271 ^ w33985;
	assign w34071 = w34082 & w34072;
	assign w34069 = w34071 ^ w34079;
	assign w34068 = w34077 & w34069;
	assign w34033 = w34068 ^ w34043;
	assign w34067 = w34033 ^ w34035;
	assign w33991 = w34068 ^ w34092;
	assign w34064 = w34033 ^ w33986;
	assign w34059 = w34073 & w47276;
	assign w34058 = w34064 & w34094;
	assign w34057 = w34067 & w34106;
	assign w34056 = w34077 & w34096;
	assign w34000 = w34056 ^ w34057;
	assign w34055 = w34065 & w34097;
	assign w34050 = w34073 & w34105;
	assign w34049 = w34064 & w34109;
	assign w34016 = w34058 ^ w34049;
	assign w34048 = w34067 & w34102;
	assign w34018 = w34056 ^ w34048;
	assign w34047 = w34077 & w34103;
	assign w34046 = w34065 & w34108;
	assign w44797 = w34057 ^ w34058;
	assign w44799 = w34071 ^ w34089;
	assign w34063 = w44799 ^ w34041;
	assign w34061 = w34063 & w34100;
	assign w44798 = w34059 ^ w34061;
	assign w34052 = w34063 & w34104;
	assign w34030 = w47275 ^ w44799;
	assign w34070 = w34030 ^ w33993;
	assign w33983 = w34030 ^ w33991;
	assign w33990 = w34020 ^ w33983;
	assign w34066 = w33987 ^ w33990;
	assign w34062 = w33983 ^ w33984;
	assign w34060 = w34070 & w34099;
	assign w34054 = w34062 & w34095;
	assign w34039 = w34054 ^ w44797;
	assign w34015 = w34054 ^ w34057;
	assign w34012 = ~w34015;
	assign w34011 = w34054 ^ w34055;
	assign w34005 = w34050 ^ w34039;
	assign w34002 = ~w34005;
	assign w33999 = w34055 ^ w34039;
	assign w34053 = w34066 & w34098;
	assign w34031 = w34049 ^ w34053;
	assign w34009 = ~w34031;
	assign w34008 = w34009 ^ w34047;
	assign w34004 = w34008 ^ w44798;
	assign w34007 = w34046 ^ w34004;
	assign w34051 = w34070 & w34101;
	assign w34045 = w34062 & w34110;
	assign w34044 = w34066 & w34107;
	assign w34010 = w34055 ^ w34044;
	assign w34006 = ~w34010;
	assign w34111 = w34006 ^ w34007;
	assign w44796 = w34045 ^ w34046;
	assign w34027 = w34051 ^ w44796;
	assign w34003 = w34027 ^ w34004;
	assign w49266 = w34002 ^ w34003;
	assign w7885 = w49266 ^ w45417;
	assign w34028 = w34052 ^ w34027;
	assign w49269 = w34028 ^ w33999;
	assign w34032 = w34060 ^ w34028;
	assign w34001 = w34059 ^ w34032;
	assign w49267 = w34000 ^ w34001;
	assign w7730 = ~w49267;
	assign w34037 = w34061 ^ w34032;
	assign w34112 = w34037 ^ w34011;
	assign w8003 = w49262 ^ w49267;
	assign w8006 = w49261 ^ w49266;
	assign w7859 = ~w8006;
	assign w7857 = w7859 ^ w49274;
	assign w7971 = w49264 ^ w49269;
	assign w7834 = w7971 ^ w45542;
	assign w7867 = ~w8003;
	assign w7729 = w7730 ^ w49261;
	assign w8058 = w7728 ^ w7729;
	assign w49268 = w44797 ^ w34037;
	assign w7999 = w49263 ^ w49268;
	assign w7732 = w49268 ^ w49262;
	assign w8057 = w7731 ^ w7732;
	assign w7841 = ~w7999;
	assign w34014 = w34018 ^ w44796;
	assign w34017 = w44798 ^ w34014;
	assign w34114 = w34016 ^ w34017;
	assign w34013 = w34009 ^ w34014;
	assign w34113 = w34012 ^ w34013;
	assign w7726 = w34113 ^ w45410;
	assign w8059 = w7725 ^ w7726;
	assign w49265 = ~w34113;
	assign w8010 = w45417 ^ w49265;
	assign w45782 = ~w34111;
	assign w7995 = w45415 ^ w45782;
	assign w7856 = w7995 ^ w45549;
	assign w7854 = ~w7856;
	assign w7863 = w7995 ^ w7989;
	assign w7883 = w45782 ^ w49263;
	assign w45783 = ~w34112;
	assign w7853 = w45783 ^ w45782;
	assign w45784 = ~w34114;
	assign w8011 = w45410 ^ w45784;
	assign w45918 = ~w7488;
	assign w7479 = w45918 ^ w45722;
	assign w49015 = w7479 ^ w7480;
	assign w7451 = w45918 ^ w45430;
	assign w49033 = w7450 ^ w7451;
	assign w47259 = w49033 ^ w45166;
	assign w7713 = w47253 ^ w47259;
	assign w7640 = w47259 ^ w47258;
	assign w7705 = w7640 ^ w7707;
	assign w7448 = w45918 ^ w49097;
	assign w7446 = w7447 ^ w7448;
	assign w49035 = ~w7446;
	assign w47257 = w49035 ^ w1495;
	assign w7623 = w47259 ^ w47257;
	assign w7625 = w47258 ^ w7623;
	assign w7704 = w7623 ^ w7712;
	assign w7701 = w47254 ^ w7625;
	assign w7698 = w47255 ^ w7625;
	assign w7703 = w47260 ^ w7704;
	assign w7696 = w7705 & w7703;
	assign w7647 = w7690 ^ w7696;
	assign w7700 = w7630 ^ w7625;
	assign w7692 = w7707 & w7700;
	assign w7694 = w7713 & w7698;
	assign w7628 = w7694 ^ w7624;
	assign w7600 = w47257 ^ w47258;
	assign w7702 = w7623 ^ w7586;
	assign w7689 = w7711 & w7702;
	assign w7691 = w7712 & w7701;
	assign w7627 = w7691 ^ w7625;
	assign w7599 = w7690 ^ w7691;
	assign w7646 = w7599 ^ w7600;
	assign w7645 = w7646 ^ w7628;
	assign w47277 = w49015 ^ w1476;
	assign w18833 = w47277 ^ w47283;
	assign w18814 = w18833 & w18818;
	assign w18831 = w47277 ^ w47282;
	assign w18832 = w47280 ^ w47277;
	assign w18811 = w18832 & w18821;
	assign w18747 = w18811 ^ w18745;
	assign w18824 = w18743 ^ w18832;
	assign w18744 = w47279 ^ w47277;
	assign w18706 = w18746 ^ w18744;
	assign w18822 = w18743 ^ w18706;
	assign w18809 = w18831 & w18822;
	assign w18827 = w18744 ^ w18750;
	assign w18812 = w18827 & w18820;
	assign w18825 = w18760 ^ w18827;
	assign w18823 = w47284 ^ w18824;
	assign w18816 = w18825 & w18823;
	assign w18748 = w18814 ^ w18744;
	assign w18828 = w18832 ^ w18760;
	assign w18817 = w18824 & w18828;
	assign w18749 = w18817 ^ w18746;
	assign w18753 = w18749 ^ w18747;
	assign w18758 = w47277 ^ w18753;
	assign w7706 = w47259 ^ w7710;
	assign w7693 = w7710 & w7706;
	assign w7687 = w7693 ^ w7645;
	assign w43792 = w7689 ^ w7695;
	assign w7639 = w43792 ^ w7624;
	assign w7685 = w7647 ^ w7639;
	assign w43793 = w7689 ^ w7692;
	assign w7642 = w7690 ^ w43793;
	assign w7598 = w7693 ^ w7642;
	assign w7680 = w47259 ^ w7598;
	assign w7602 = w7628 ^ w43793;
	assign w7686 = w7602 ^ w7627;
	assign w44154 = w18809 ^ w18815;
	assign w18721 = w18753 ^ w44154;
	assign w18764 = w47279 ^ w18721;
	assign w18759 = w44154 ^ w18744;
	assign w7708 = w7712 ^ w7640;
	assign w7697 = w7704 & w7708;
	assign w7629 = w7697 ^ w7626;
	assign w7633 = w7629 ^ w7627;
	assign w7638 = w47253 ^ w7633;
	assign w7688 = w7647 ^ w7638;
	assign w7684 = w7688 & w7687;
	assign w7683 = w7684 ^ w7686;
	assign w7682 = w7685 & w7683;
	assign w7590 = w7682 ^ w7638;
	assign w7593 = w7682 ^ w7694;
	assign w7589 = w7593 ^ w7629;
	assign w7588 = w47255 ^ w7589;
	assign w7601 = w7633 ^ w43792;
	assign w7644 = w47255 ^ w7601;
	assign w7679 = w7684 ^ w7644;
	assign w7678 = w7679 & w7680;
	assign w7676 = w7684 ^ w7678;
	assign w7675 = w7686 & w7676;
	assign w7673 = w7675 ^ w7683;
	assign w7677 = w7678 ^ w7686;
	assign w7663 = w7677 & w47260;
	assign w7681 = w7682 ^ w7644;
	assign w7672 = w7681 & w7673;
	assign w7596 = w7678 ^ w7695;
	assign w7591 = w7596 ^ w7692;
	assign w7595 = w7672 ^ w7696;
	assign w7660 = w7681 & w7700;
	assign w7654 = w7677 & w7709;
	assign w7651 = w7681 & w7707;
	assign w7637 = w7672 ^ w7647;
	assign w7668 = w7637 ^ w7590;
	assign w7671 = w7637 ^ w7639;
	assign w7662 = w7668 & w7698;
	assign w7661 = w7671 & w7710;
	assign w7604 = w7660 ^ w7661;
	assign w7653 = w7668 & w7713;
	assign w7620 = w7662 ^ w7653;
	assign w7652 = w7671 & w7706;
	assign w7622 = w7660 ^ w7652;
	assign w7597 = w7678 ^ w7642;
	assign w43795 = w7661 ^ w7662;
	assign w43797 = w7675 ^ w7693;
	assign w7667 = w43797 ^ w7645;
	assign w7665 = w7667 & w7704;
	assign w43796 = w7663 ^ w7665;
	assign w7656 = w7667 & w7708;
	assign w7634 = w47259 ^ w43797;
	assign w7674 = w7634 ^ w7597;
	assign w7664 = w7674 & w7703;
	assign w7655 = w7674 & w7705;
	assign w7587 = w7634 ^ w7595;
	assign w7666 = w7587 ^ w7588;
	assign w7649 = w7666 & w7714;
	assign w7658 = w7666 & w7699;
	assign w7643 = w7658 ^ w43795;
	assign w7619 = w7658 ^ w7661;
	assign w7616 = ~w7619;
	assign w7609 = w7654 ^ w7643;
	assign w7606 = ~w7609;
	assign w7594 = w7624 ^ w7587;
	assign w7670 = w7591 ^ w7594;
	assign w7648 = w7670 & w7711;
	assign w7657 = w7670 & w7702;
	assign w7635 = w7653 ^ w7657;
	assign w7613 = ~w7635;
	assign w7612 = w7613 ^ w7651;
	assign w7608 = w7612 ^ w43796;
	assign w7592 = w47253 ^ w7589;
	assign w7669 = w7591 ^ w7592;
	assign w7659 = w7669 & w7701;
	assign w7615 = w7658 ^ w7659;
	assign w7614 = w7659 ^ w7648;
	assign w7610 = ~w7614;
	assign w7603 = w7659 ^ w7643;
	assign w7650 = w7669 & w7712;
	assign w7611 = w7650 ^ w7608;
	assign w7715 = w7610 ^ w7611;
	assign w43794 = w7649 ^ w7650;
	assign w7631 = w7655 ^ w43794;
	assign w7607 = w7631 ^ w7608;
	assign w49310 = w7606 ^ w7607;
	assign w7632 = w7656 ^ w7631;
	assign w7636 = w7664 ^ w7632;
	assign w7641 = w7665 ^ w7636;
	assign w7716 = w7641 ^ w7615;
	assign w49312 = w43795 ^ w7641;
	assign w7605 = w7663 ^ w7636;
	assign w49311 = w7604 ^ w7605;
	assign w7736 = w49311 ^ w49310;
	assign w49313 = w7632 ^ w7603;
	assign w7967 = w49309 ^ w49313;
	assign w7774 = w7967 ^ w49311;
	assign w8039 = w7774 ^ w7775;
	assign w7984 = w49308 ^ w49312;
	assign w7924 = w7992 ^ w7984;
	assign w7985 = w49306 ^ w49310;
	assign w7926 = w7987 ^ w7985;
	assign w7939 = w7982 ^ w49312;
	assign w7618 = w7622 ^ w43794;
	assign w7621 = w43796 ^ w7618;
	assign w7718 = w7620 ^ w7621;
	assign w7617 = w7613 ^ w7618;
	assign w7717 = w7616 ^ w7617;
	assign w45197 = ~w7716;
	assign w7990 = w45630 ^ w45197;
	assign w7945 = w7990 ^ w45264;
	assign w45198 = ~w7717;
	assign w7719 = w7982 ^ w45198;
	assign w8062 = w7719 ^ w7720;
	assign w7777 = w45198 ^ w49302;
	assign w7997 = w45631 ^ w45198;
	assign w45199 = ~w7718;
	assign w7734 = w45199 ^ w45258;
	assign w8017 = w45632 ^ w45199;
	assign w45200 = ~w7715;
	assign w7961 = w7963 ^ w45200;
	assign w18819 = w18744 ^ w18834;
	assign w18810 = w18834 & w18819;
	assign w18719 = w18810 ^ w18811;
	assign w18766 = w18719 ^ w18720;
	assign w18767 = w18810 ^ w18816;
	assign w18808 = w18767 ^ w18758;
	assign w18805 = w18767 ^ w18759;
	assign w18765 = w18766 ^ w18748;
	assign w18807 = w18813 ^ w18765;
	assign w18804 = w18808 & w18807;
	assign w18799 = w18804 ^ w18764;
	assign w44155 = w18809 ^ w18812;
	assign w18722 = w18748 ^ w44155;
	assign w18806 = w18722 ^ w18747;
	assign w18803 = w18804 ^ w18806;
	assign w18802 = w18805 & w18803;
	assign w18801 = w18802 ^ w18764;
	assign w18780 = w18801 & w18820;
	assign w18771 = w18801 & w18827;
	assign w18710 = w18802 ^ w18758;
	assign w18713 = w18802 ^ w18814;
	assign w18709 = w18713 ^ w18749;
	assign w18712 = w47277 ^ w18709;
	assign w18708 = w47279 ^ w18709;
	assign w18762 = w18810 ^ w44155;
	assign w18718 = w18813 ^ w18762;
	assign w18800 = w47283 ^ w18718;
	assign w18798 = w18799 & w18800;
	assign w18717 = w18798 ^ w18762;
	assign w18716 = w18798 ^ w18815;
	assign w18711 = w18716 ^ w18812;
	assign w18789 = w18711 ^ w18712;
	assign w18779 = w18789 & w18821;
	assign w18770 = w18789 & w18832;
	assign w18796 = w18804 ^ w18798;
	assign w18795 = w18806 & w18796;
	assign w18793 = w18795 ^ w18803;
	assign w18792 = w18801 & w18793;
	assign w18715 = w18792 ^ w18816;
	assign w18797 = w18798 ^ w18806;
	assign w18783 = w18797 & w47284;
	assign w18774 = w18797 & w18829;
	assign w44159 = w18795 ^ w18813;
	assign w18787 = w44159 ^ w18765;
	assign w18785 = w18787 & w18824;
	assign w44158 = w18783 ^ w18785;
	assign w18776 = w18787 & w18828;
	assign w18757 = w18792 ^ w18767;
	assign w18788 = w18757 ^ w18710;
	assign w18773 = w18788 & w18833;
	assign w18782 = w18788 & w18818;
	assign w18791 = w18757 ^ w18759;
	assign w18781 = w18791 & w18830;
	assign w18772 = w18791 & w18826;
	assign w18742 = w18780 ^ w18772;
	assign w18724 = w18780 ^ w18781;
	assign w18740 = w18782 ^ w18773;
	assign w44157 = w18781 ^ w18782;
	assign w18754 = w47283 ^ w44159;
	assign w18794 = w18754 ^ w18717;
	assign w18775 = w18794 & w18825;
	assign w18784 = w18794 & w18823;
	assign w18707 = w18754 ^ w18715;
	assign w18786 = w18707 ^ w18708;
	assign w18714 = w18744 ^ w18707;
	assign w18778 = w18786 & w18819;
	assign w18769 = w18786 & w18834;
	assign w18735 = w18778 ^ w18779;
	assign w44156 = w18769 ^ w18770;
	assign w18751 = w18775 ^ w44156;
	assign w18738 = w18742 ^ w44156;
	assign w18741 = w44158 ^ w18738;
	assign w18790 = w18711 ^ w18714;
	assign w18768 = w18790 & w18831;
	assign w18777 = w18790 & w18822;
	assign w18734 = w18779 ^ w18768;
	assign w18730 = ~w18734;
	assign w18755 = w18773 ^ w18777;
	assign w18733 = ~w18755;
	assign w18737 = w18733 ^ w18738;
	assign w18732 = w18733 ^ w18771;
	assign w18728 = w18732 ^ w44158;
	assign w18727 = w18751 ^ w18728;
	assign w18838 = w18740 ^ w18741;
	assign w45406 = ~w18838;
	assign w18739 = w18778 ^ w18781;
	assign w18736 = ~w18739;
	assign w18837 = w18736 ^ w18737;
	assign w45413 = ~w18837;
	assign w18763 = w18778 ^ w44157;
	assign w18723 = w18779 ^ w18763;
	assign w18729 = w18774 ^ w18763;
	assign w18726 = ~w18729;
	assign w49278 = w18726 ^ w18727;
	assign w18731 = w18770 ^ w18728;
	assign w18835 = w18730 ^ w18731;
	assign w45411 = ~w18835;
	assign w18752 = w18776 ^ w18751;
	assign w49281 = w18752 ^ w18723;
	assign w18756 = w18784 ^ w18752;
	assign w18761 = w18785 ^ w18756;
	assign w18836 = w18761 ^ w18735;
	assign w7977 = w49281 ^ w49296;
	assign w7750 = w7977 ^ w49294;
	assign w7746 = ~w7977;
	assign w7747 = w7746 ^ w49293;
	assign w7744 = w7746 ^ w45715;
	assign w7833 = w8031 ^ w7977;
	assign w49280 = w44157 ^ w18761;
	assign w18725 = w18783 ^ w18756;
	assign w49279 = w18724 ^ w18725;
	assign w45412 = ~w18836;
	assign w45919 = ~w7495;
	assign w7283 = w45919 ^ w45268;
	assign w7565 = w7283 ^ w7284;
	assign w48921 = w7565 ^ w7557;
	assign w7419 = w45919 ^ w49059;
	assign w48935 = w7419 ^ w7420;
	assign w47357 = w48935 ^ w1587;
	assign w19146 = w47359 ^ w47357;
	assign w19221 = w19146 ^ w19236;
	assign w19234 = w47360 ^ w47357;
	assign w19226 = w19145 ^ w19234;
	assign w19225 = w47364 ^ w19226;
	assign w19230 = w19234 ^ w19162;
	assign w19229 = w19146 ^ w19152;
	assign w19227 = w19162 ^ w19229;
	assign w19235 = w47357 ^ w47363;
	assign w19233 = w47357 ^ w47362;
	assign w19216 = w19235 & w19220;
	assign w19150 = w19216 ^ w19146;
	assign w19108 = w19148 ^ w19146;
	assign w19212 = w19236 & w19221;
	assign w19219 = w19226 & w19230;
	assign w19151 = w19219 ^ w19148;
	assign w19213 = w19234 & w19223;
	assign w19149 = w19213 ^ w19147;
	assign w19155 = w19151 ^ w19149;
	assign w19160 = w47357 ^ w19155;
	assign w19218 = w19227 & w19225;
	assign w19169 = w19212 ^ w19218;
	assign w19210 = w19169 ^ w19160;
	assign w19121 = w19212 ^ w19213;
	assign w19168 = w19121 ^ w19122;
	assign w19167 = w19168 ^ w19150;
	assign w19209 = w19215 ^ w19167;
	assign w7440 = w45919 ^ w49042;
	assign w48924 = w7439 ^ w7440;
	assign w47371 = w48921 ^ w1573;
	assign w33751 = w47371 ^ w47369;
	assign w33753 = w47370 ^ w33751;
	assign w33829 = w47366 ^ w33753;
	assign w33826 = w47367 ^ w33753;
	assign w33828 = w33758 ^ w33753;
	assign w33834 = w47371 ^ w33838;
	assign w33768 = w47371 ^ w47370;
	assign w33833 = w33768 ^ w33835;
	assign w33841 = w47365 ^ w47371;
	assign w33822 = w33841 & w33826;
	assign w33756 = w33822 ^ w33752;
	assign w33821 = w33838 & w33834;
	assign w33820 = w33835 & w33828;
	assign w47368 = w48924 ^ w1576;
	assign w33754 = w47368 ^ w47366;
	assign w33840 = w47368 ^ w47365;
	assign w33836 = w33840 ^ w33768;
	assign w33832 = w33751 ^ w33840;
	assign w33831 = w47372 ^ w33832;
	assign w33842 = w47370 ^ w47368;
	assign w33827 = w33752 ^ w33842;
	assign w33714 = w33754 ^ w33752;
	assign w33830 = w33751 ^ w33714;
	assign w33713 = w33754 ^ w47367;
	assign w33837 = w47372 ^ w33713;
	assign w33825 = w33832 & w33836;
	assign w33757 = w33825 ^ w33754;
	assign w33824 = w33833 & w33831;
	assign w33823 = w47372 & w33837;
	assign w33819 = w33840 & w33829;
	assign w33755 = w33819 ^ w33753;
	assign w33761 = w33757 ^ w33755;
	assign w33766 = w47365 ^ w33761;
	assign w33818 = w33842 & w33827;
	assign w33775 = w33818 ^ w33824;
	assign w33816 = w33775 ^ w33766;
	assign w33727 = w33818 ^ w33819;
	assign w33774 = w33727 ^ w33728;
	assign w33773 = w33774 ^ w33756;
	assign w33815 = w33821 ^ w33773;
	assign w33817 = w33839 & w33830;
	assign w33812 = w33816 & w33815;
	assign w19214 = w19229 & w19222;
	assign w19206 = w19210 & w19209;
	assign w44782 = w33817 ^ w33823;
	assign w33729 = w33761 ^ w44782;
	assign w33772 = w47367 ^ w33729;
	assign w33807 = w33812 ^ w33772;
	assign w33767 = w44782 ^ w33752;
	assign w33813 = w33775 ^ w33767;
	assign w44783 = w33817 ^ w33820;
	assign w33770 = w33818 ^ w44783;
	assign w33726 = w33821 ^ w33770;
	assign w33808 = w47371 ^ w33726;
	assign w33806 = w33807 & w33808;
	assign w33724 = w33806 ^ w33823;
	assign w33719 = w33724 ^ w33820;
	assign w33804 = w33812 ^ w33806;
	assign w33725 = w33806 ^ w33770;
	assign w33730 = w33756 ^ w44783;
	assign w33814 = w33730 ^ w33755;
	assign w33805 = w33806 ^ w33814;
	assign w33811 = w33812 ^ w33814;
	assign w33810 = w33813 & w33811;
	assign w33809 = w33810 ^ w33772;
	assign w33721 = w33810 ^ w33822;
	assign w33717 = w33721 ^ w33757;
	assign w33720 = w47365 ^ w33717;
	assign w33797 = w33719 ^ w33720;
	assign w33718 = w33810 ^ w33766;
	assign w33716 = w47367 ^ w33717;
	assign w33803 = w33814 & w33804;
	assign w33801 = w33803 ^ w33811;
	assign w33800 = w33809 & w33801;
	assign w33765 = w33800 ^ w33775;
	assign w33799 = w33765 ^ w33767;
	assign w33723 = w33800 ^ w33824;
	assign w33796 = w33765 ^ w33718;
	assign w33791 = w33805 & w47372;
	assign w33790 = w33796 & w33826;
	assign w33789 = w33799 & w33838;
	assign w33788 = w33809 & w33828;
	assign w33732 = w33788 ^ w33789;
	assign w33787 = w33797 & w33829;
	assign w33782 = w33805 & w33837;
	assign w33781 = w33796 & w33841;
	assign w33748 = w33790 ^ w33781;
	assign w33780 = w33799 & w33834;
	assign w33750 = w33788 ^ w33780;
	assign w33779 = w33809 & w33835;
	assign w33778 = w33797 & w33840;
	assign w44785 = w33789 ^ w33790;
	assign w44787 = w33803 ^ w33821;
	assign w33795 = w44787 ^ w33773;
	assign w33793 = w33795 & w33832;
	assign w44786 = w33791 ^ w33793;
	assign w33784 = w33795 & w33836;
	assign w33762 = w47371 ^ w44787;
	assign w33802 = w33762 ^ w33725;
	assign w33715 = w33762 ^ w33723;
	assign w33722 = w33752 ^ w33715;
	assign w33798 = w33719 ^ w33722;
	assign w33794 = w33715 ^ w33716;
	assign w33792 = w33802 & w33831;
	assign w33786 = w33794 & w33827;
	assign w33771 = w33786 ^ w44785;
	assign w33747 = w33786 ^ w33789;
	assign w33744 = ~w33747;
	assign w33743 = w33786 ^ w33787;
	assign w33737 = w33782 ^ w33771;
	assign w33734 = ~w33737;
	assign w33731 = w33787 ^ w33771;
	assign w33785 = w33798 & w33830;
	assign w33763 = w33781 ^ w33785;
	assign w33741 = ~w33763;
	assign w33740 = w33741 ^ w33779;
	assign w33736 = w33740 ^ w44786;
	assign w33739 = w33778 ^ w33736;
	assign w33783 = w33802 & w33833;
	assign w33777 = w33794 & w33842;
	assign w33776 = w33798 & w33839;
	assign w33742 = w33787 ^ w33776;
	assign w33738 = ~w33742;
	assign w33843 = w33738 ^ w33739;
	assign w7797 = w45419 ^ w33843;
	assign w7828 = w33843 ^ w49280;
	assign w49182 = w7827 ^ w7828;
	assign w47183 = w49182 ^ w1633;
	assign w49286 = ~w33843;
	assign w8005 = w45411 ^ w49286;
	assign w7781 = w8005 ^ w8000;
	assign w49206 = w45419 ^ w7781;
	assign w7799 = w8005 ^ w45720;
	assign w7808 = w8005 ^ w7983;
	assign w49191 = w45412 ^ w7808;
	assign w47159 = w49206 ^ w1657;
	assign w47174 = w49191 ^ w1642;
	assign w44784 = w33777 ^ w33778;
	assign w33759 = w33783 ^ w44784;
	assign w33760 = w33784 ^ w33759;
	assign w49288 = w33760 ^ w33731;
	assign w7820 = w49288 ^ w45412;
	assign w49184 = w7819 ^ w7820;
	assign w47181 = w49184 ^ w1635;
	assign w33764 = w33792 ^ w33760;
	assign w33733 = w33791 ^ w33764;
	assign w49284 = w33732 ^ w33733;
	assign w7749 = ~w49284;
	assign w7748 = w7749 ^ w49278;
	assign w8050 = w7747 ^ w7748;
	assign w33769 = w33793 ^ w33764;
	assign w49285 = w44785 ^ w33769;
	assign w7751 = w49285 ^ w49279;
	assign w8049 = w7750 ^ w7751;
	assign w7800 = w49291 ^ w49285;
	assign w33844 = w33769 ^ w33743;
	assign w49287 = ~w33844;
	assign w7976 = w49288 ^ w49292;
	assign w7752 = w7976 ^ w45714;
	assign w7757 = ~w7976;
	assign w7754 = w7757 ^ w49294;
	assign w7758 = w7757 ^ w49295;
	assign w7998 = w45412 ^ w49287;
	assign w7780 = w7998 ^ w7994;
	assign w49207 = w45420 ^ w7780;
	assign w7798 = w7998 ^ w45721;
	assign w7796 = ~w7798;
	assign w7807 = w7998 ^ w7969;
	assign w49192 = w49281 ^ w7807;
	assign w49199 = w7796 ^ w7797;
	assign w47158 = w49207 ^ w1658;
	assign w8012 = w49280 ^ w49285;
	assign w7784 = ~w8012;
	assign w7782 = w7784 ^ w8009;
	assign w7809 = w8012 ^ w7994;
	assign w49190 = w45411 ^ w7809;
	assign w7823 = w33844 ^ w45411;
	assign w7821 = w7822 ^ w7823;
	assign w49183 = ~w7821;
	assign w47182 = w49183 ^ w1634;
	assign w7795 = w45420 ^ w33844;
	assign w49198 = w7799 ^ w7800;
	assign w33735 = w33759 ^ w33736;
	assign w49283 = w33734 ^ w33735;
	assign w8027 = w49278 ^ w49283;
	assign w7803 = ~w8027;
	assign w7801 = w7803 ^ w49293;
	assign w7812 = w7803 ^ w8009;
	assign w7788 = w8027 ^ w8023;
	assign w49203 = w49289 ^ w7788;
	assign w8020 = w49279 ^ w49284;
	assign w7787 = ~w8020;
	assign w7810 = w7787 ^ w8000;
	assign w7785 = w7787 ^ w8019;
	assign w49181 = w8049 ^ w8000;
	assign w47184 = w49181 ^ w1632;
	assign w18430 = w47184 ^ w47181;
	assign w18344 = w47184 ^ w47182;
	assign w18303 = w18344 ^ w47183;
	assign w7972 = w49281 ^ w49288;
	assign w7818 = w8031 ^ w7972;
	assign w7779 = w7983 ^ w7972;
	assign w49208 = w49292 ^ w7779;
	assign w47157 = w49208 ^ w1659;
	assign w30804 = w47159 ^ w47157;
	assign w49180 = w8050 ^ w8009;
	assign w47185 = w49180 ^ w1631;
	assign w7756 = ~w49283;
	assign w7831 = w7756 ^ w45413;
	assign w49179 = w7830 ^ w7831;
	assign w47186 = w49179 ^ w1630;
	assign w18318 = w47185 ^ w47186;
	assign w18432 = w47186 ^ w47184;
	assign w47173 = w49192 ^ w1643;
	assign w47175 = w49190 ^ w1641;
	assign w33618 = w47175 ^ w47173;
	assign w7759 = w49290 ^ w7749;
	assign w8046 = w7758 ^ w7759;
	assign w49197 = w8046 ^ w8012;
	assign w47162 = w49203 ^ w1654;
	assign w30891 = w47157 ^ w47162;
	assign w47166 = w49199 ^ w1650;
	assign w47167 = w49198 ^ w1649;
	assign w47168 = w49197 ^ w1648;
	assign w18210 = w47168 ^ w47166;
	assign w18169 = w18210 ^ w47167;
	assign w49185 = w45406 ^ w7818;
	assign w47180 = w49185 ^ w1636;
	assign w33624 = w47180 ^ w47174;
	assign w33701 = w33618 ^ w33624;
	assign w33704 = w47175 ^ w33624;
	assign w18342 = w47183 ^ w47181;
	assign w18417 = w18342 ^ w18432;
	assign w18408 = w18432 & w18417;
	assign w7755 = w49289 ^ w7756;
	assign w8047 = w7754 ^ w7755;
	assign w49196 = w8047 ^ w8020;
	assign w47169 = w49196 ^ w1647;
	assign w33746 = w33750 ^ w44784;
	assign w33749 = w44786 ^ w33746;
	assign w33846 = w33748 ^ w33749;
	assign w33745 = w33741 ^ w33746;
	assign w33845 = w33744 ^ w33745;
	assign w7745 = w33845 ^ w45406;
	assign w8051 = w7744 ^ w7745;
	assign w7802 = w45421 ^ w33845;
	assign w49195 = w7801 ^ w7802;
	assign w49282 = ~w33845;
	assign w49178 = w8051 ^ w8023;
	assign w47187 = w49178 ^ w1629;
	assign w18358 = w47187 ^ w47186;
	assign w18426 = w18430 ^ w18358;
	assign w8034 = w45413 ^ w49282;
	assign w7814 = w8034 ^ w8019;
	assign w49187 = w49278 ^ w7814;
	assign w7792 = w8034 ^ w8031;
	assign w7790 = ~w7792;
	assign w47178 = w49187 ^ w1638;
	assign w33705 = w47173 ^ w47178;
	assign w18341 = w47187 ^ w47185;
	assign w18343 = w47186 ^ w18341;
	assign w18419 = w47182 ^ w18343;
	assign w18416 = w47183 ^ w18343;
	assign w18409 = w18430 & w18419;
	assign w18345 = w18409 ^ w18343;
	assign w18317 = w18408 ^ w18409;
	assign w18422 = w18341 ^ w18430;
	assign w18415 = w18422 & w18426;
	assign w18347 = w18415 ^ w18344;
	assign w18351 = w18347 ^ w18345;
	assign w18356 = w47181 ^ w18351;
	assign w47170 = w49195 ^ w1646;
	assign w18298 = w47170 ^ w47168;
	assign w18184 = w47169 ^ w47170;
	assign w18364 = w18317 ^ w18318;
	assign w18304 = w18344 ^ w18342;
	assign w18420 = w18341 ^ w18304;
	assign w19224 = w19145 ^ w19108;
	assign w19211 = w19233 & w19224;
	assign w44171 = w19211 ^ w19214;
	assign w19124 = w19150 ^ w44171;
	assign w19208 = w19124 ^ w19149;
	assign w19205 = w19206 ^ w19208;
	assign w19164 = w19212 ^ w44171;
	assign w19120 = w19215 ^ w19164;
	assign w19202 = w47363 ^ w19120;
	assign w44174 = w19211 ^ w19217;
	assign w19123 = w19155 ^ w44174;
	assign w19166 = w47359 ^ w19123;
	assign w19201 = w19206 ^ w19166;
	assign w19161 = w44174 ^ w19146;
	assign w19207 = w19169 ^ w19161;
	assign w18431 = w47181 ^ w47187;
	assign w18412 = w18431 & w18416;
	assign w18346 = w18412 ^ w18342;
	assign w18363 = w18364 ^ w18346;
	assign w19204 = w19207 & w19205;
	assign w19203 = w19204 ^ w19166;
	assign w19112 = w19204 ^ w19160;
	assign w19115 = w19204 ^ w19216;
	assign w19111 = w19115 ^ w19151;
	assign w19114 = w47357 ^ w19111;
	assign w19173 = w19203 & w19229;
	assign w19182 = w19203 & w19222;
	assign w19110 = w47359 ^ w19111;
	assign w19200 = w19201 & w19202;
	assign w19118 = w19200 ^ w19217;
	assign w19113 = w19118 ^ w19214;
	assign w19119 = w19200 ^ w19164;
	assign w19198 = w19206 ^ w19200;
	assign w19197 = w19208 & w19198;
	assign w19195 = w19197 ^ w19205;
	assign w19194 = w19203 & w19195;
	assign w19159 = w19194 ^ w19169;
	assign w19193 = w19159 ^ w19161;
	assign w19191 = w19113 ^ w19114;
	assign w19190 = w19159 ^ w19112;
	assign w19184 = w19190 & w19220;
	assign w19172 = w19191 & w19234;
	assign w44173 = w19197 ^ w19215;
	assign w19189 = w44173 ^ w19167;
	assign w19187 = w19189 & w19226;
	assign w19178 = w19189 & w19230;
	assign w19156 = w47363 ^ w44173;
	assign w19196 = w19156 ^ w19119;
	assign w19177 = w19196 & w19227;
	assign w19199 = w19200 ^ w19208;
	assign w19176 = w19199 & w19231;
	assign w19186 = w19196 & w19225;
	assign w19117 = w19194 ^ w19218;
	assign w19109 = w19156 ^ w19117;
	assign w19188 = w19109 ^ w19110;
	assign w19180 = w19188 & w19221;
	assign w19171 = w19188 & w19236;
	assign w44172 = w19171 ^ w19172;
	assign w19153 = w19177 ^ w44172;
	assign w19154 = w19178 ^ w19153;
	assign w19158 = w19186 ^ w19154;
	assign w19163 = w19187 ^ w19158;
	assign w19116 = w19146 ^ w19109;
	assign w19192 = w19113 ^ w19116;
	assign w19170 = w19192 & w19233;
	assign w18429 = w47181 ^ w47186;
	assign w18407 = w18429 & w18420;
	assign w19185 = w19199 & w47364;
	assign w19127 = w19185 ^ w19158;
	assign w44176 = w19185 ^ w19187;
	assign w19183 = w19193 & w19232;
	assign w19126 = w19182 ^ w19183;
	assign w49271 = w19126 ^ w19127;
	assign w7742 = w49271 ^ w7730;
	assign w7996 = w49271 ^ w49275;
	assign w7868 = w7859 ^ w7996;
	assign w49148 = w8058 ^ w7996;
	assign w47217 = w49148 ^ w1663;
	assign w7838 = w7841 ^ w7996;
	assign w19141 = w19180 ^ w19183;
	assign w19138 = ~w19141;
	assign w44175 = w19183 ^ w19184;
	assign w49272 = w44175 ^ w19163;
	assign w7840 = ~w49272;
	assign w7855 = w7840 ^ w49268;
	assign w7991 = w49272 ^ w49276;
	assign w49149 = w8057 ^ w7991;
	assign w47216 = w49149 ^ w1664;
	assign w7837 = w7995 ^ w7991;
	assign w7865 = w7867 ^ w7991;
	assign w19165 = w19180 ^ w44175;
	assign w19131 = w19176 ^ w19165;
	assign w19128 = ~w19131;
	assign w49166 = w7854 ^ w7855;
	assign w47199 = w49166 ^ w1681;
	assign w19181 = w19191 & w19223;
	assign w19137 = w19180 ^ w19181;
	assign w19125 = w19181 ^ w19165;
	assign w19238 = w19163 ^ w19137;
	assign w19136 = w19181 ^ w19170;
	assign w49273 = w19154 ^ w19125;
	assign w19132 = ~w19136;
	assign w7970 = w49273 ^ w49277;
	assign w7839 = w7970 ^ w7840;
	assign w49173 = w7838 ^ w7839;
	assign w7861 = w7970 ^ w45783;
	assign w7850 = w8011 ^ w7970;
	assign w7978 = w49269 ^ w49273;
	assign w7739 = w7978 ^ w49275;
	assign w7737 = w7978 ^ w45543;
	assign w7743 = ~w7978;
	assign w7741 = w7743 ^ w49276;
	assign w8052 = w7741 ^ w7742;
	assign w7860 = w8011 ^ w7978;
	assign w49161 = w45544 ^ w7860;
	assign w47204 = w49161 ^ w1676;
	assign w49165 = w8052 ^ w7999;
	assign w47192 = w49173 ^ w1688;
	assign w49160 = w7861 ^ w7862;
	assign w47205 = w49160 ^ w1675;
	assign w7846 = w7970 ^ w49271;
	assign w47200 = w49165 ^ w1680;
	assign w7879 = w7989 ^ w7970;
	assign w49152 = w49269 ^ w7879;
	assign w47213 = w49152 ^ w1667;
	assign w18564 = w47216 ^ w47213;
	assign w45424 = ~w19238;
	assign w7835 = w49273 ^ w45424;
	assign w49176 = w7834 ^ w7835;
	assign w49159 = w45424 ^ w7863;
	assign w47206 = w49159 ^ w1674;
	assign w7988 = w45783 ^ w45424;
	assign w7880 = w7988 ^ w45542;
	assign w7851 = w7988 ^ w7971;
	assign w49168 = w49277 ^ w7851;
	assign w47189 = w49176 ^ w1691;
	assign w31026 = w47192 ^ w47189;
	assign w49151 = w7880 ^ w7881;
	assign w47214 = w49151 ^ w1666;
	assign w18478 = w47216 ^ w47214;
	assign w47197 = w49168 ^ w1683;
	assign w27856 = w47199 ^ w47197;
	assign w27944 = w47200 ^ w47197;
	assign w19179 = w19192 & w19224;
	assign w45778 = ~w33846;
	assign w7753 = w45414 ^ w45778;
	assign w8048 = w7752 ^ w7753;
	assign w49177 = w45778 ^ w7833;
	assign w47188 = w49177 ^ w1628;
	assign w18348 = w47188 ^ w47182;
	assign w18425 = w18342 ^ w18348;
	assign w18428 = w47183 ^ w18348;
	assign w18423 = w18358 ^ w18425;
	assign w18421 = w47188 ^ w18422;
	assign w18418 = w18348 ^ w18343;
	assign w18410 = w18425 & w18418;
	assign w18414 = w18423 & w18421;
	assign w18365 = w18408 ^ w18414;
	assign w18406 = w18365 ^ w18356;
	assign w49194 = w8048 ^ w8034;
	assign w8035 = w45406 ^ w45778;
	assign w7804 = w8035 ^ w7976;
	assign w49193 = w45715 ^ w7804;
	assign w7793 = w8035 ^ w7969;
	assign w49201 = w45414 ^ w7793;
	assign w47172 = w49193 ^ w1644;
	assign w18293 = w47172 ^ w18169;
	assign w18279 = w47172 & w18293;
	assign w18214 = w47172 ^ w47166;
	assign w18294 = w47167 ^ w18214;
	assign w47164 = w49201 ^ w1652;
	assign w30810 = w47164 ^ w47158;
	assign w30887 = w30804 ^ w30810;
	assign w30890 = w47159 ^ w30810;
	assign w7816 = w8035 ^ w8023;
	assign w18424 = w47187 ^ w18428;
	assign w18411 = w18428 & w18424;
	assign w18405 = w18411 ^ w18363;
	assign w18402 = w18406 & w18405;
	assign w47171 = w49194 ^ w1645;
	assign w18224 = w47171 ^ w47170;
	assign w18207 = w47171 ^ w47169;
	assign w18209 = w47170 ^ w18207;
	assign w18285 = w47166 ^ w18209;
	assign w18282 = w47167 ^ w18209;
	assign w18290 = w47171 ^ w18294;
	assign w18277 = w18294 & w18290;
	assign w18284 = w18214 ^ w18209;
	assign w44138 = w18407 ^ w18410;
	assign w18360 = w18408 ^ w44138;
	assign w18316 = w18411 ^ w18360;
	assign w18398 = w47187 ^ w18316;
	assign w18320 = w18346 ^ w44138;
	assign w18404 = w18320 ^ w18345;
	assign w18401 = w18402 ^ w18404;
	assign w18427 = w47188 ^ w18303;
	assign w18413 = w47188 & w18427;
	assign w44137 = w18407 ^ w18413;
	assign w18319 = w18351 ^ w44137;
	assign w18362 = w47183 ^ w18319;
	assign w18397 = w18402 ^ w18362;
	assign w18396 = w18397 & w18398;
	assign w18315 = w18396 ^ w18360;
	assign w18314 = w18396 ^ w18413;
	assign w18394 = w18402 ^ w18396;
	assign w18393 = w18404 & w18394;
	assign w18391 = w18393 ^ w18401;
	assign w18395 = w18396 ^ w18404;
	assign w18372 = w18395 & w18427;
	assign w18381 = w18395 & w47188;
	assign w18357 = w44137 ^ w18342;
	assign w18403 = w18365 ^ w18357;
	assign w18400 = w18403 & w18401;
	assign w18311 = w18400 ^ w18412;
	assign w18308 = w18400 ^ w18356;
	assign w18399 = w18400 ^ w18362;
	assign w18378 = w18399 & w18418;
	assign w18390 = w18399 & w18391;
	assign w18355 = w18390 ^ w18365;
	assign w18313 = w18390 ^ w18414;
	assign w18389 = w18355 ^ w18357;
	assign w18379 = w18389 & w18428;
	assign w18322 = w18378 ^ w18379;
	assign w18370 = w18389 & w18424;
	assign w18340 = w18378 ^ w18370;
	assign w18369 = w18399 & w18425;
	assign w44141 = w18393 ^ w18411;
	assign w18385 = w44141 ^ w18363;
	assign w18374 = w18385 & w18426;
	assign w18383 = w18385 & w18422;
	assign w44140 = w18381 ^ w18383;
	assign w18352 = w47187 ^ w44141;
	assign w18392 = w18352 ^ w18315;
	assign w18373 = w18392 & w18423;
	assign w18305 = w18352 ^ w18313;
	assign w18382 = w18392 & w18421;
	assign w18309 = w18314 ^ w18410;
	assign w18307 = w18311 ^ w18347;
	assign w18310 = w47181 ^ w18307;
	assign w18387 = w18309 ^ w18310;
	assign w18368 = w18387 & w18430;
	assign w18377 = w18387 & w18419;
	assign w18312 = w18342 ^ w18305;
	assign w18388 = w18309 ^ w18312;
	assign w18366 = w18388 & w18429;
	assign w18332 = w18377 ^ w18366;
	assign w18328 = ~w18332;
	assign w18375 = w18388 & w18420;
	assign w18386 = w18355 ^ w18308;
	assign w18371 = w18386 & w18431;
	assign w18353 = w18371 ^ w18375;
	assign w18331 = ~w18353;
	assign w18330 = w18331 ^ w18369;
	assign w18326 = w18330 ^ w44140;
	assign w18329 = w18368 ^ w18326;
	assign w18433 = w18328 ^ w18329;
	assign w18306 = w47183 ^ w18307;
	assign w45398 = ~w18433;
	assign w18384 = w18305 ^ w18306;
	assign w18367 = w18384 & w18432;
	assign w43550 = w18367 ^ w18368;
	assign w18336 = w18340 ^ w43550;
	assign w18339 = w44140 ^ w18336;
	assign w18335 = w18331 ^ w18336;
	assign w18349 = w18373 ^ w43550;
	assign w18325 = w18349 ^ w18326;
	assign w18350 = w18374 ^ w18349;
	assign w18354 = w18382 ^ w18350;
	assign w18359 = w18383 ^ w18354;
	assign w18323 = w18381 ^ w18354;
	assign w49463 = w18322 ^ w18323;
	assign w18376 = w18384 & w18417;
	assign w18337 = w18376 ^ w18379;
	assign w18334 = ~w18337;
	assign w18435 = w18334 ^ w18335;
	assign w18333 = w18376 ^ w18377;
	assign w18434 = w18359 ^ w18333;
	assign w45399 = ~w18434;
	assign w45400 = ~w18435;
	assign w18380 = w18386 & w18416;
	assign w18338 = w18380 ^ w18371;
	assign w18436 = w18338 ^ w18339;
	assign w44139 = w18379 ^ w18380;
	assign w18361 = w18376 ^ w44139;
	assign w18327 = w18372 ^ w18361;
	assign w18321 = w18377 ^ w18361;
	assign w49465 = w18350 ^ w18321;
	assign w8340 = w49465 ^ w45399;
	assign w18324 = ~w18327;
	assign w49462 = w18324 ^ w18325;
	assign w49464 = w44139 ^ w18359;
	assign w45401 = ~w18436;
	assign w19175 = w19190 & w19235;
	assign w19142 = w19184 ^ w19175;
	assign w19157 = w19175 ^ w19179;
	assign w19135 = ~w19157;
	assign w19134 = w19135 ^ w19173;
	assign w19130 = w19134 ^ w44176;
	assign w19133 = w19172 ^ w19130;
	assign w19237 = w19132 ^ w19133;
	assign w19129 = w19153 ^ w19130;
	assign w49270 = w19128 ^ w19129;
	assign w7740 = w49270 ^ w49266;
	assign w8053 = w7739 ^ w7740;
	assign w49164 = w8053 ^ w8003;
	assign w8001 = w49270 ^ w49274;
	assign w7870 = w8010 ^ w8001;
	assign w49155 = w49261 ^ w7870;
	assign w47210 = w49155 ^ w1670;
	assign w12801 = w47205 ^ w47210;
	assign w7845 = w8003 ^ w8001;
	assign w49172 = w7845 ^ w7846;
	assign w47193 = w49172 ^ w1687;
	assign w47201 = w49164 ^ w1679;
	assign w7884 = w8001 ^ w45543;
	assign w49147 = w7884 ^ w7885;
	assign w47218 = w49147 ^ w1662;
	assign w18566 = w47218 ^ w47216;
	assign w18563 = w47213 ^ w47218;
	assign w18452 = w47217 ^ w47218;
	assign w45423 = ~w19237;
	assign w49174 = w45423 ^ w7837;
	assign w7986 = w45423 ^ w45549;
	assign w7882 = w7986 ^ w49276;
	assign w7836 = w7988 ^ w7986;
	assign w49175 = w45416 ^ w7836;
	assign w7852 = w7989 ^ w45423;
	assign w49167 = w7852 ^ w7853;
	assign w49150 = w7882 ^ w7883;
	assign w47215 = w49150 ^ w1665;
	assign w47190 = w49175 ^ w1690;
	assign w30940 = w47192 ^ w47190;
	assign w47191 = w49174 ^ w1689;
	assign w30938 = w47191 ^ w47189;
	assign w30900 = w30940 ^ w30938;
	assign w30899 = w30940 ^ w47191;
	assign w7864 = w7999 ^ w7986;
	assign w47198 = w49167 ^ w1682;
	assign w27858 = w47200 ^ w47198;
	assign w27862 = w47204 ^ w47198;
	assign w27939 = w27856 ^ w27862;
	assign w27942 = w47199 ^ w27862;
	assign w27818 = w27858 ^ w27856;
	assign w27817 = w27858 ^ w47199;
	assign w27941 = w47204 ^ w27817;
	assign w27927 = w47204 & w27941;
	assign w49158 = w45415 ^ w7864;
	assign w47207 = w49158 ^ w1673;
	assign w12714 = w47207 ^ w47205;
	assign w18476 = w47215 ^ w47213;
	assign w18438 = w18478 ^ w18476;
	assign w18551 = w18476 ^ w18566;
	assign w18542 = w18566 & w18551;
	assign w18437 = w18478 ^ w47215;
	assign w45892 = ~w7972;
	assign w7811 = w45892 ^ w49280;
	assign w7794 = w45892 ^ w49296;
	assign w7813 = w45892 ^ w49279;
	assign w49188 = w7812 ^ w7813;
	assign w49200 = w7794 ^ w7795;
	assign w49189 = w7810 ^ w7811;
	assign w47177 = w49188 ^ w1639;
	assign w33594 = w47177 ^ w47178;
	assign w47176 = w49189 ^ w1640;
	assign w33620 = w47176 ^ w47174;
	assign w33706 = w47176 ^ w47173;
	assign w33708 = w47178 ^ w47176;
	assign w33693 = w33618 ^ w33708;
	assign w33580 = w33620 ^ w33618;
	assign w33579 = w33620 ^ w47175;
	assign w33703 = w47180 ^ w33579;
	assign w33689 = w47180 & w33703;
	assign w33684 = w33708 & w33693;
	assign w7817 = w45892 ^ w45413;
	assign w47165 = w49200 ^ w1651;
	assign w18208 = w47167 ^ w47165;
	assign w18170 = w18210 ^ w18208;
	assign w18286 = w18207 ^ w18170;
	assign w18296 = w47168 ^ w47165;
	assign w18275 = w18296 & w18285;
	assign w18211 = w18275 ^ w18209;
	assign w18283 = w18208 ^ w18298;
	assign w18274 = w18298 & w18283;
	assign w18295 = w47165 ^ w47170;
	assign w18273 = w18295 & w18286;
	assign w18288 = w18207 ^ w18296;
	assign w18287 = w47172 ^ w18288;
	assign w18297 = w47165 ^ w47171;
	assign w18278 = w18297 & w18282;
	assign w18212 = w18278 ^ w18208;
	assign w18291 = w18208 ^ w18214;
	assign w18289 = w18224 ^ w18291;
	assign w18280 = w18289 & w18287;
	assign w18276 = w18291 & w18284;
	assign w18292 = w18296 ^ w18224;
	assign w18281 = w18288 & w18292;
	assign w18213 = w18281 ^ w18210;
	assign w7815 = w7816 ^ w7817;
	assign w49186 = ~w7815;
	assign w47179 = w49186 ^ w1637;
	assign w33617 = w47179 ^ w47177;
	assign w33619 = w47178 ^ w33617;
	assign w33695 = w47174 ^ w33619;
	assign w33692 = w47175 ^ w33619;
	assign w33694 = w33624 ^ w33619;
	assign w33700 = w47179 ^ w33704;
	assign w33698 = w33617 ^ w33706;
	assign w33697 = w47180 ^ w33698;
	assign w33634 = w47179 ^ w47178;
	assign w33699 = w33634 ^ w33701;
	assign w33702 = w33706 ^ w33634;
	assign w33696 = w33617 ^ w33580;
	assign w33707 = w47173 ^ w47179;
	assign w33691 = w33698 & w33702;
	assign w33623 = w33691 ^ w33620;
	assign w33690 = w33699 & w33697;
	assign w33641 = w33684 ^ w33690;
	assign w33688 = w33707 & w33692;
	assign w33622 = w33688 ^ w33618;
	assign w33687 = w33704 & w33700;
	assign w33686 = w33701 & w33694;
	assign w33685 = w33706 & w33695;
	assign w33621 = w33685 ^ w33619;
	assign w33627 = w33623 ^ w33621;
	assign w33632 = w47173 ^ w33627;
	assign w33682 = w33641 ^ w33632;
	assign w33593 = w33684 ^ w33685;
	assign w33640 = w33593 ^ w33594;
	assign w33639 = w33640 ^ w33622;
	assign w33681 = w33687 ^ w33639;
	assign w33683 = w33705 & w33696;
	assign w33678 = w33682 & w33681;
	assign w44131 = w18273 ^ w18276;
	assign w18186 = w18212 ^ w44131;
	assign w18270 = w18186 ^ w18211;
	assign w18226 = w18274 ^ w44131;
	assign w18182 = w18277 ^ w18226;
	assign w18264 = w47171 ^ w18182;
	assign w44134 = w18273 ^ w18279;
	assign w18223 = w44134 ^ w18208;
	assign w18231 = w18274 ^ w18280;
	assign w18269 = w18231 ^ w18223;
	assign w18217 = w18213 ^ w18211;
	assign w18222 = w47165 ^ w18217;
	assign w18272 = w18231 ^ w18222;
	assign w18185 = w18217 ^ w44134;
	assign w18228 = w47167 ^ w18185;
	assign w44777 = w33683 ^ w33689;
	assign w33633 = w44777 ^ w33618;
	assign w33679 = w33641 ^ w33633;
	assign w33595 = w33627 ^ w44777;
	assign w33638 = w47175 ^ w33595;
	assign w33673 = w33678 ^ w33638;
	assign w44778 = w33683 ^ w33686;
	assign w33636 = w33684 ^ w44778;
	assign w33592 = w33687 ^ w33636;
	assign w33674 = w47179 ^ w33592;
	assign w33672 = w33673 & w33674;
	assign w33591 = w33672 ^ w33636;
	assign w33590 = w33672 ^ w33689;
	assign w33585 = w33590 ^ w33686;
	assign w33670 = w33678 ^ w33672;
	assign w33596 = w33622 ^ w44778;
	assign w33680 = w33596 ^ w33621;
	assign w33671 = w33672 ^ w33680;
	assign w33677 = w33678 ^ w33680;
	assign w33676 = w33679 & w33677;
	assign w33675 = w33676 ^ w33638;
	assign w33587 = w33676 ^ w33688;
	assign w33583 = w33587 ^ w33623;
	assign w33586 = w47173 ^ w33583;
	assign w33663 = w33585 ^ w33586;
	assign w33584 = w33676 ^ w33632;
	assign w33582 = w47175 ^ w33583;
	assign w33669 = w33680 & w33670;
	assign w33667 = w33669 ^ w33677;
	assign w33666 = w33675 & w33667;
	assign w33631 = w33666 ^ w33641;
	assign w33665 = w33631 ^ w33633;
	assign w33589 = w33666 ^ w33690;
	assign w33662 = w33631 ^ w33584;
	assign w33657 = w33671 & w47180;
	assign w33656 = w33662 & w33692;
	assign w33655 = w33665 & w33704;
	assign w33654 = w33675 & w33694;
	assign w33598 = w33654 ^ w33655;
	assign w33653 = w33663 & w33695;
	assign w33648 = w33671 & w33703;
	assign w33647 = w33662 & w33707;
	assign w33614 = w33656 ^ w33647;
	assign w33646 = w33665 & w33700;
	assign w33616 = w33654 ^ w33646;
	assign w33645 = w33675 & w33701;
	assign w33644 = w33663 & w33706;
	assign w44779 = w33655 ^ w33656;
	assign w44781 = w33669 ^ w33687;
	assign w33628 = w47179 ^ w44781;
	assign w33668 = w33628 ^ w33591;
	assign w33649 = w33668 & w33699;
	assign w33658 = w33668 & w33697;
	assign w33581 = w33628 ^ w33589;
	assign w33588 = w33618 ^ w33581;
	assign w33664 = w33585 ^ w33588;
	assign w33651 = w33664 & w33696;
	assign w33629 = w33647 ^ w33651;
	assign w33607 = ~w33629;
	assign w33606 = w33607 ^ w33645;
	assign w33660 = w33581 ^ w33582;
	assign w33643 = w33660 & w33708;
	assign w33642 = w33664 & w33705;
	assign w33608 = w33653 ^ w33642;
	assign w33604 = ~w33608;
	assign w43594 = w33643 ^ w33644;
	assign w33625 = w33649 ^ w43594;
	assign w33612 = w33616 ^ w43594;
	assign w33611 = w33607 ^ w33612;
	assign w33652 = w33660 & w33693;
	assign w33609 = w33652 ^ w33653;
	assign w33637 = w33652 ^ w44779;
	assign w33603 = w33648 ^ w33637;
	assign w33600 = ~w33603;
	assign w33597 = w33653 ^ w33637;
	assign w33613 = w33652 ^ w33655;
	assign w33610 = ~w33613;
	assign w33711 = w33610 ^ w33611;
	assign w33661 = w44781 ^ w33639;
	assign w33659 = w33661 & w33698;
	assign w33650 = w33661 & w33702;
	assign w33626 = w33650 ^ w33625;
	assign w33630 = w33658 ^ w33626;
	assign w33635 = w33659 ^ w33630;
	assign w49448 = w44779 ^ w33635;
	assign w33710 = w33635 ^ w33609;
	assign w33599 = w33657 ^ w33630;
	assign w49447 = w33598 ^ w33599;
	assign w49451 = w33626 ^ w33597;
	assign w49450 = ~w33710;
	assign w44780 = w33657 ^ w33659;
	assign w33615 = w44780 ^ w33612;
	assign w33712 = w33614 ^ w33615;
	assign w33602 = w33606 ^ w44780;
	assign w33605 = w33644 ^ w33602;
	assign w33709 = w33604 ^ w33605;
	assign w33601 = w33625 ^ w33602;
	assign w49446 = w33600 ^ w33601;
	assign w49449 = ~w33709;
	assign w18183 = w18274 ^ w18275;
	assign w18230 = w18183 ^ w18184;
	assign w18229 = w18230 ^ w18212;
	assign w18271 = w18277 ^ w18229;
	assign w18268 = w18272 & w18271;
	assign w18263 = w18268 ^ w18228;
	assign w18267 = w18268 ^ w18270;
	assign w18266 = w18269 & w18267;
	assign w18265 = w18266 ^ w18228;
	assign w18244 = w18265 & w18284;
	assign w18177 = w18266 ^ w18278;
	assign w18174 = w18266 ^ w18222;
	assign w18235 = w18265 & w18291;
	assign w18262 = w18263 & w18264;
	assign w18260 = w18268 ^ w18262;
	assign w18259 = w18270 & w18260;
	assign w18181 = w18262 ^ w18226;
	assign w18257 = w18259 ^ w18267;
	assign w18256 = w18265 & w18257;
	assign w18221 = w18256 ^ w18231;
	assign w18252 = w18221 ^ w18174;
	assign w18246 = w18252 & w18282;
	assign w18255 = w18221 ^ w18223;
	assign w18245 = w18255 & w18294;
	assign w18188 = w18244 ^ w18245;
	assign w18237 = w18252 & w18297;
	assign w18204 = w18246 ^ w18237;
	assign w18236 = w18255 & w18290;
	assign w18206 = w18244 ^ w18236;
	assign w18261 = w18262 ^ w18270;
	assign w18238 = w18261 & w18293;
	assign w18247 = w18261 & w47172;
	assign w44133 = w18259 ^ w18277;
	assign w18218 = w47171 ^ w44133;
	assign w18258 = w18218 ^ w18181;
	assign w18239 = w18258 & w18289;
	assign w18248 = w18258 & w18287;
	assign w44135 = w18245 ^ w18246;
	assign w18251 = w44133 ^ w18229;
	assign w18249 = w18251 & w18288;
	assign w44136 = w18247 ^ w18249;
	assign w18180 = w18262 ^ w18279;
	assign w18175 = w18180 ^ w18276;
	assign w18179 = w18256 ^ w18280;
	assign w18171 = w18218 ^ w18179;
	assign w18178 = w18208 ^ w18171;
	assign w18254 = w18175 ^ w18178;
	assign w18232 = w18254 & w18295;
	assign w18241 = w18254 & w18286;
	assign w18219 = w18237 ^ w18241;
	assign w18197 = ~w18219;
	assign w18196 = w18197 ^ w18235;
	assign w18192 = w18196 ^ w44136;
	assign w18173 = w18177 ^ w18213;
	assign w18172 = w47167 ^ w18173;
	assign w18250 = w18171 ^ w18172;
	assign w18233 = w18250 & w18298;
	assign w18242 = w18250 & w18283;
	assign w18203 = w18242 ^ w18245;
	assign w18200 = ~w18203;
	assign w18227 = w18242 ^ w44135;
	assign w18193 = w18238 ^ w18227;
	assign w18190 = ~w18193;
	assign w18240 = w18251 & w18292;
	assign w18176 = w47165 ^ w18173;
	assign w18253 = w18175 ^ w18176;
	assign w18234 = w18253 & w18296;
	assign w44132 = w18233 ^ w18234;
	assign w18215 = w18239 ^ w44132;
	assign w18216 = w18240 ^ w18215;
	assign w18220 = w18248 ^ w18216;
	assign w18225 = w18249 ^ w18220;
	assign w49509 = w44135 ^ w18225;
	assign w18189 = w18247 ^ w18220;
	assign w49508 = w18188 ^ w18189;
	assign w8253 = w49509 ^ w49508;
	assign w18191 = w18215 ^ w18192;
	assign w49507 = w18190 ^ w18191;
	assign w18202 = w18206 ^ w44132;
	assign w18205 = w44136 ^ w18202;
	assign w18302 = w18204 ^ w18205;
	assign w18201 = w18197 ^ w18202;
	assign w18243 = w18253 & w18285;
	assign w18199 = w18242 ^ w18243;
	assign w18198 = w18243 ^ w18232;
	assign w18300 = w18225 ^ w18199;
	assign w18194 = ~w18198;
	assign w18187 = w18243 ^ w18227;
	assign w49510 = w18216 ^ w18187;
	assign w18301 = w18200 ^ w18201;
	assign w18195 = w18234 ^ w18192;
	assign w18299 = w18194 ^ w18195;
	assign w45394 = ~w18299;
	assign w45395 = ~w18300;
	assign w8401 = w45395 ^ w45394;
	assign w45396 = ~w18301;
	assign w45397 = ~w18302;
	assign w45779 = ~w33711;
	assign w45780 = ~w33712;
	assign w19174 = w19193 & w19228;
	assign w19144 = w19182 ^ w19174;
	assign w19140 = w19144 ^ w44172;
	assign w19139 = w19135 ^ w19140;
	assign w19143 = w44176 ^ w19140;
	assign w19240 = w19142 ^ w19143;
	assign w19239 = w19138 ^ w19139;
	assign w45418 = ~w19240;
	assign w7738 = w45418 ^ w45784;
	assign w8054 = w7737 ^ w7738;
	assign w49169 = w45418 ^ w7850;
	assign w47196 = w49169 ^ w1684;
	assign w30944 = w47196 ^ w47190;
	assign w31021 = w30938 ^ w30944;
	assign w31024 = w47191 ^ w30944;
	assign w31023 = w47196 ^ w30899;
	assign w31009 = w47196 & w31023;
	assign w8008 = w45418 ^ w45544;
	assign w49162 = w8054 ^ w8010;
	assign w7848 = w8010 ^ w8008;
	assign w47203 = w49162 ^ w1677;
	assign w27855 = w47203 ^ w47201;
	assign w27938 = w47203 ^ w27942;
	assign w27936 = w27855 ^ w27944;
	assign w27935 = w47204 ^ w27936;
	assign w27934 = w27855 ^ w27818;
	assign w27945 = w47197 ^ w47203;
	assign w27925 = w27942 & w27938;
	assign w7874 = w8008 ^ w7971;
	assign w49153 = w45410 ^ w7874;
	assign w47212 = w49153 ^ w1668;
	assign w7886 = w8008 ^ w7980;
	assign w49145 = w45784 ^ w7886;
	assign w47220 = w49145 ^ w1660;
	assign w18482 = w47220 ^ w47214;
	assign w18562 = w47215 ^ w18482;
	assign w18561 = w47220 ^ w18437;
	assign w18559 = w18476 ^ w18482;
	assign w12720 = w47212 ^ w47206;
	assign w12797 = w12714 ^ w12720;
	assign w12800 = w47207 ^ w12720;
	assign w18547 = w47220 & w18561;
	assign w45425 = ~w19239;
	assign w7858 = w45425 ^ w34113;
	assign w7849 = w7970 ^ w45425;
	assign w49170 = w7848 ^ w7849;
	assign w8004 = w45425 ^ w45543;
	assign w49146 = w8059 ^ w8004;
	assign w47219 = w49146 ^ w1661;
	assign w18492 = w47219 ^ w47218;
	assign w18565 = w47213 ^ w47219;
	assign w18558 = w47219 ^ w18562;
	assign w18545 = w18562 & w18558;
	assign w18560 = w18564 ^ w18492;
	assign w49163 = w7857 ^ w7858;
	assign w47202 = w49163 ^ w1678;
	assign w27857 = w47202 ^ w27855;
	assign w27933 = w47198 ^ w27857;
	assign w27930 = w47199 ^ w27857;
	assign w27932 = w27862 ^ w27857;
	assign w27872 = w47203 ^ w47202;
	assign w27937 = w27872 ^ w27939;
	assign w27940 = w27944 ^ w27872;
	assign w27946 = w47202 ^ w47200;
	assign w27931 = w27856 ^ w27946;
	assign w27832 = w47201 ^ w47202;
	assign w27943 = w47197 ^ w47202;
	assign w27929 = w27936 & w27940;
	assign w27861 = w27929 ^ w27858;
	assign w27928 = w27937 & w27935;
	assign w27926 = w27945 & w27930;
	assign w27860 = w27926 ^ w27856;
	assign w27924 = w27939 & w27932;
	assign w27923 = w27944 & w27933;
	assign w27859 = w27923 ^ w27857;
	assign w27865 = w27861 ^ w27859;
	assign w27870 = w47197 ^ w27865;
	assign w27922 = w27946 & w27931;
	assign w27879 = w27922 ^ w27928;
	assign w27920 = w27879 ^ w27870;
	assign w27831 = w27922 ^ w27923;
	assign w27878 = w27831 ^ w27832;
	assign w27877 = w27878 ^ w27860;
	assign w27919 = w27925 ^ w27877;
	assign w27921 = w27943 & w27934;
	assign w27916 = w27920 & w27919;
	assign w18475 = w47219 ^ w47217;
	assign w18477 = w47218 ^ w18475;
	assign w18550 = w47215 ^ w18477;
	assign w18554 = w18475 ^ w18438;
	assign w18556 = w18475 ^ w18564;
	assign w18555 = w47220 ^ w18556;
	assign w18552 = w18482 ^ w18477;
	assign w18544 = w18559 & w18552;
	assign w18553 = w47214 ^ w18477;
	assign w18543 = w18564 & w18553;
	assign w18479 = w18543 ^ w18477;
	assign w18546 = w18565 & w18550;
	assign w18480 = w18546 ^ w18476;
	assign w18541 = w18563 & w18554;
	assign w18549 = w18556 & w18560;
	assign w18481 = w18549 ^ w18478;
	assign w18485 = w18481 ^ w18479;
	assign w47195 = w49170 ^ w1685;
	assign w30937 = w47195 ^ w47193;
	assign w31020 = w47195 ^ w31024;
	assign w31018 = w30937 ^ w31026;
	assign w31017 = w47196 ^ w31018;
	assign w31016 = w30937 ^ w30900;
	assign w31027 = w47189 ^ w47195;
	assign w31007 = w31024 & w31020;
	assign w7847 = w8006 ^ w8004;
	assign w18451 = w18542 ^ w18543;
	assign w18498 = w18451 ^ w18452;
	assign w18497 = w18498 ^ w18480;
	assign w18539 = w18545 ^ w18497;
	assign w49171 = w49270 ^ w7847;
	assign w47194 = w49171 ^ w1686;
	assign w30939 = w47194 ^ w30937;
	assign w31015 = w47190 ^ w30939;
	assign w31012 = w47191 ^ w30939;
	assign w31014 = w30944 ^ w30939;
	assign w30954 = w47195 ^ w47194;
	assign w31019 = w30954 ^ w31021;
	assign w31022 = w31026 ^ w30954;
	assign w31028 = w47194 ^ w47192;
	assign w31013 = w30938 ^ w31028;
	assign w30914 = w47193 ^ w47194;
	assign w31025 = w47189 ^ w47194;
	assign w31011 = w31018 & w31022;
	assign w30943 = w31011 ^ w30940;
	assign w31010 = w31019 & w31017;
	assign w31008 = w31027 & w31012;
	assign w30942 = w31008 ^ w30938;
	assign w31006 = w31021 & w31014;
	assign w31005 = w31026 & w31015;
	assign w30941 = w31005 ^ w30939;
	assign w30947 = w30943 ^ w30941;
	assign w30952 = w47189 ^ w30947;
	assign w31004 = w31028 & w31013;
	assign w30961 = w31004 ^ w31010;
	assign w31002 = w30961 ^ w30952;
	assign w30913 = w31004 ^ w31005;
	assign w30960 = w30913 ^ w30914;
	assign w30959 = w30960 ^ w30942;
	assign w31001 = w31007 ^ w30959;
	assign w31003 = w31025 & w31016;
	assign w30998 = w31002 & w31001;
	assign w44142 = w18541 ^ w18547;
	assign w18453 = w18485 ^ w44142;
	assign w18496 = w47215 ^ w18453;
	assign w18491 = w44142 ^ w18476;
	assign w44143 = w18541 ^ w18544;
	assign w18494 = w18542 ^ w44143;
	assign w18454 = w18480 ^ w44143;
	assign w18538 = w18454 ^ w18479;
	assign w44534 = w27921 ^ w27924;
	assign w27834 = w27860 ^ w44534;
	assign w27918 = w27834 ^ w27859;
	assign w27915 = w27916 ^ w27918;
	assign w27874 = w27922 ^ w44534;
	assign w27830 = w27925 ^ w27874;
	assign w27912 = w47203 ^ w27830;
	assign w44537 = w27921 ^ w27927;
	assign w27833 = w27865 ^ w44537;
	assign w27876 = w47199 ^ w27833;
	assign w27911 = w27916 ^ w27876;
	assign w27910 = w27911 & w27912;
	assign w27909 = w27910 ^ w27918;
	assign w27908 = w27916 ^ w27910;
	assign w27829 = w27910 ^ w27874;
	assign w27828 = w27910 ^ w27927;
	assign w27823 = w27828 ^ w27924;
	assign w27907 = w27918 & w27908;
	assign w27905 = w27907 ^ w27915;
	assign w27895 = w27909 & w47204;
	assign w27886 = w27909 & w27941;
	assign w44536 = w27907 ^ w27925;
	assign w27899 = w44536 ^ w27877;
	assign w27897 = w27899 & w27936;
	assign w27888 = w27899 & w27940;
	assign w27866 = w47203 ^ w44536;
	assign w27906 = w27866 ^ w27829;
	assign w27896 = w27906 & w27935;
	assign w27887 = w27906 & w27937;
	assign w27871 = w44537 ^ w27856;
	assign w27917 = w27879 ^ w27871;
	assign w27914 = w27917 & w27915;
	assign w27913 = w27914 ^ w27876;
	assign w27825 = w27914 ^ w27926;
	assign w27821 = w27825 ^ w27861;
	assign w27824 = w47197 ^ w27821;
	assign w27901 = w27823 ^ w27824;
	assign w27822 = w27914 ^ w27870;
	assign w27820 = w47199 ^ w27821;
	assign w27904 = w27913 & w27905;
	assign w27869 = w27904 ^ w27879;
	assign w27903 = w27869 ^ w27871;
	assign w27827 = w27904 ^ w27928;
	assign w27819 = w27866 ^ w27827;
	assign w27826 = w27856 ^ w27819;
	assign w27902 = w27823 ^ w27826;
	assign w27900 = w27869 ^ w27822;
	assign w27898 = w27819 ^ w27820;
	assign w27894 = w27900 & w27930;
	assign w27893 = w27903 & w27942;
	assign w27892 = w27913 & w27932;
	assign w27836 = w27892 ^ w27893;
	assign w27891 = w27901 & w27933;
	assign w27890 = w27898 & w27931;
	assign w27851 = w27890 ^ w27893;
	assign w27848 = ~w27851;
	assign w27847 = w27890 ^ w27891;
	assign w27889 = w27902 & w27934;
	assign w27885 = w27900 & w27945;
	assign w27867 = w27885 ^ w27889;
	assign w27852 = w27894 ^ w27885;
	assign w27845 = ~w27867;
	assign w27884 = w27903 & w27938;
	assign w27854 = w27892 ^ w27884;
	assign w27883 = w27913 & w27939;
	assign w27844 = w27845 ^ w27883;
	assign w27882 = w27901 & w27944;
	assign w27881 = w27898 & w27946;
	assign w27880 = w27902 & w27943;
	assign w27846 = w27891 ^ w27880;
	assign w27842 = ~w27846;
	assign w44535 = w27881 ^ w27882;
	assign w27863 = w27887 ^ w44535;
	assign w27864 = w27888 ^ w27863;
	assign w27868 = w27896 ^ w27864;
	assign w27873 = w27897 ^ w27868;
	assign w27948 = w27873 ^ w27847;
	assign w27837 = w27895 ^ w27868;
	assign w49491 = w27836 ^ w27837;
	assign w27850 = w27854 ^ w44535;
	assign w27849 = w27845 ^ w27850;
	assign w27949 = w27848 ^ w27849;
	assign w44538 = w27893 ^ w27894;
	assign w49492 = w44538 ^ w27873;
	assign w27875 = w27890 ^ w44538;
	assign w27841 = w27886 ^ w27875;
	assign w27838 = ~w27841;
	assign w27835 = w27891 ^ w27875;
	assign w49493 = w27864 ^ w27835;
	assign w44539 = w27895 ^ w27897;
	assign w27853 = w44539 ^ w27850;
	assign w27950 = w27852 ^ w27853;
	assign w27840 = w27844 ^ w44539;
	assign w27843 = w27882 ^ w27840;
	assign w27947 = w27842 ^ w27843;
	assign w27839 = w27863 ^ w27840;
	assign w49490 = w27838 ^ w27839;
	assign w44666 = w31003 ^ w31009;
	assign w30953 = w44666 ^ w30938;
	assign w30999 = w30961 ^ w30953;
	assign w30915 = w30947 ^ w44666;
	assign w30958 = w47191 ^ w30915;
	assign w30993 = w30998 ^ w30958;
	assign w44667 = w31003 ^ w31006;
	assign w30956 = w31004 ^ w44667;
	assign w30912 = w31007 ^ w30956;
	assign w30994 = w47195 ^ w30912;
	assign w30992 = w30993 & w30994;
	assign w30911 = w30992 ^ w30956;
	assign w30910 = w30992 ^ w31009;
	assign w30905 = w30910 ^ w31006;
	assign w30990 = w30998 ^ w30992;
	assign w30916 = w30942 ^ w44667;
	assign w31000 = w30916 ^ w30941;
	assign w30991 = w30992 ^ w31000;
	assign w30997 = w30998 ^ w31000;
	assign w30996 = w30999 & w30997;
	assign w30995 = w30996 ^ w30958;
	assign w30907 = w30996 ^ w31008;
	assign w30903 = w30907 ^ w30943;
	assign w30906 = w47189 ^ w30903;
	assign w30983 = w30905 ^ w30906;
	assign w30904 = w30996 ^ w30952;
	assign w30902 = w47191 ^ w30903;
	assign w30989 = w31000 & w30990;
	assign w30987 = w30989 ^ w30997;
	assign w30986 = w30995 & w30987;
	assign w30951 = w30986 ^ w30961;
	assign w30985 = w30951 ^ w30953;
	assign w30909 = w30986 ^ w31010;
	assign w30982 = w30951 ^ w30904;
	assign w30977 = w30991 & w47196;
	assign w30976 = w30982 & w31012;
	assign w30975 = w30985 & w31024;
	assign w30974 = w30995 & w31014;
	assign w30918 = w30974 ^ w30975;
	assign w30973 = w30983 & w31015;
	assign w30968 = w30991 & w31023;
	assign w30967 = w30982 & w31027;
	assign w30934 = w30976 ^ w30967;
	assign w30966 = w30985 & w31020;
	assign w30936 = w30974 ^ w30966;
	assign w30965 = w30995 & w31021;
	assign w30964 = w30983 & w31026;
	assign w44668 = w30975 ^ w30976;
	assign w44670 = w30989 ^ w31007;
	assign w30948 = w47195 ^ w44670;
	assign w30988 = w30948 ^ w30911;
	assign w30969 = w30988 & w31019;
	assign w30978 = w30988 & w31017;
	assign w30901 = w30948 ^ w30909;
	assign w30908 = w30938 ^ w30901;
	assign w30984 = w30905 ^ w30908;
	assign w30971 = w30984 & w31016;
	assign w30949 = w30967 ^ w30971;
	assign w30927 = ~w30949;
	assign w30926 = w30927 ^ w30965;
	assign w30980 = w30901 ^ w30902;
	assign w30963 = w30980 & w31028;
	assign w30962 = w30984 & w31025;
	assign w30928 = w30973 ^ w30962;
	assign w30924 = ~w30928;
	assign w43585 = w30963 ^ w30964;
	assign w30932 = w30936 ^ w43585;
	assign w30931 = w30927 ^ w30932;
	assign w30945 = w30969 ^ w43585;
	assign w30972 = w30980 & w31013;
	assign w30929 = w30972 ^ w30973;
	assign w30957 = w30972 ^ w44668;
	assign w30923 = w30968 ^ w30957;
	assign w30920 = ~w30923;
	assign w30917 = w30973 ^ w30957;
	assign w30933 = w30972 ^ w30975;
	assign w30930 = ~w30933;
	assign w31031 = w30930 ^ w30931;
	assign w30981 = w44670 ^ w30959;
	assign w30979 = w30981 & w31018;
	assign w30970 = w30981 & w31022;
	assign w30946 = w30970 ^ w30945;
	assign w30950 = w30978 ^ w30946;
	assign w30955 = w30979 ^ w30950;
	assign w49477 = w44668 ^ w30955;
	assign w31030 = w30955 ^ w30929;
	assign w30919 = w30977 ^ w30950;
	assign w49476 = w30918 ^ w30919;
	assign w49478 = w30946 ^ w30917;
	assign w8458 = w49465 ^ w49478;
	assign w8205 = ~w8458;
	assign w8209 = w8458 ^ w49476;
	assign w44669 = w30977 ^ w30979;
	assign w30935 = w44669 ^ w30932;
	assign w31032 = w30934 ^ w30935;
	assign w30922 = w30926 ^ w44669;
	assign w30925 = w30964 ^ w30922;
	assign w31029 = w30924 ^ w30925;
	assign w30921 = w30945 ^ w30922;
	assign w49475 = w30920 ^ w30921;
	assign w8206 = w8205 ^ w49475;
	assign w18557 = w18492 ^ w18559;
	assign w18548 = w18557 & w18555;
	assign w18499 = w18542 ^ w18548;
	assign w18537 = w18499 ^ w18491;
	assign w7872 = w8011 ^ w8004;
	assign w18490 = w47213 ^ w18485;
	assign w18540 = w18499 ^ w18490;
	assign w18536 = w18540 & w18539;
	assign w18531 = w18536 ^ w18496;
	assign w18535 = w18536 ^ w18538;
	assign w18534 = w18537 & w18535;
	assign w18445 = w18534 ^ w18546;
	assign w18441 = w18445 ^ w18481;
	assign w18444 = w47213 ^ w18441;
	assign w18442 = w18534 ^ w18490;
	assign w18533 = w18534 ^ w18496;
	assign w18503 = w18533 & w18559;
	assign w18512 = w18533 & w18552;
	assign w18440 = w47215 ^ w18441;
	assign w18450 = w18545 ^ w18494;
	assign w18532 = w47219 ^ w18450;
	assign w18530 = w18531 & w18532;
	assign w18448 = w18530 ^ w18547;
	assign w18443 = w18448 ^ w18544;
	assign w18521 = w18443 ^ w18444;
	assign w18449 = w18530 ^ w18494;
	assign w18502 = w18521 & w18564;
	assign w18511 = w18521 & w18553;
	assign w18529 = w18530 ^ w18538;
	assign w18515 = w18529 & w47220;
	assign w18506 = w18529 & w18561;
	assign w18528 = w18536 ^ w18530;
	assign w18527 = w18538 & w18528;
	assign w18525 = w18527 ^ w18535;
	assign w18524 = w18533 & w18525;
	assign w18489 = w18524 ^ w18499;
	assign w18447 = w18524 ^ w18548;
	assign w18523 = w18489 ^ w18491;
	assign w18513 = w18523 & w18562;
	assign w18504 = w18523 & w18558;
	assign w18474 = w18512 ^ w18504;
	assign w18456 = w18512 ^ w18513;
	assign w44147 = w18527 ^ w18545;
	assign w18519 = w44147 ^ w18497;
	assign w18517 = w18519 & w18556;
	assign w44146 = w18515 ^ w18517;
	assign w18508 = w18519 & w18560;
	assign w18486 = w47219 ^ w44147;
	assign w18439 = w18486 ^ w18447;
	assign w18526 = w18486 ^ w18449;
	assign w18507 = w18526 & w18557;
	assign w18516 = w18526 & w18555;
	assign w18518 = w18439 ^ w18440;
	assign w18501 = w18518 & w18566;
	assign w18510 = w18518 & w18551;
	assign w18471 = w18510 ^ w18513;
	assign w18468 = ~w18471;
	assign w18467 = w18510 ^ w18511;
	assign w18446 = w18476 ^ w18439;
	assign w18522 = w18443 ^ w18446;
	assign w18500 = w18522 & w18563;
	assign w18466 = w18511 ^ w18500;
	assign w18462 = ~w18466;
	assign w18509 = w18522 & w18554;
	assign w44144 = w18501 ^ w18502;
	assign w18483 = w18507 ^ w44144;
	assign w18470 = w18474 ^ w44144;
	assign w18473 = w44146 ^ w18470;
	assign w18520 = w18489 ^ w18442;
	assign w18514 = w18520 & w18550;
	assign w18505 = w18520 & w18565;
	assign w18472 = w18514 ^ w18505;
	assign w18570 = w18472 ^ w18473;
	assign w18487 = w18505 ^ w18509;
	assign w18465 = ~w18487;
	assign w18464 = w18465 ^ w18503;
	assign w18460 = w18464 ^ w44146;
	assign w18463 = w18502 ^ w18460;
	assign w18567 = w18462 ^ w18463;
	assign w18469 = w18465 ^ w18470;
	assign w18569 = w18468 ^ w18469;
	assign w44145 = w18513 ^ w18514;
	assign w18495 = w18510 ^ w44145;
	assign w18461 = w18506 ^ w18495;
	assign w18458 = ~w18461;
	assign w18455 = w18511 ^ w18495;
	assign w45402 = ~w18567;
	assign w8504 = w45402 ^ w49449;
	assign w45404 = ~w18569;
	assign w45405 = ~w18570;
	assign w18484 = w18508 ^ w18483;
	assign w49445 = w18484 ^ w18455;
	assign w8452 = w49445 ^ w49451;
	assign w18488 = w18516 ^ w18484;
	assign w18457 = w18515 ^ w18488;
	assign w49443 = w18456 ^ w18457;
	assign w8516 = w49443 ^ w49447;
	assign w18493 = w18517 ^ w18488;
	assign w49444 = w44145 ^ w18493;
	assign w8507 = w49444 ^ w49448;
	assign w18568 = w18493 ^ w18467;
	assign w8242 = w8452 ^ w49443;
	assign w8398 = ~w8516;
	assign w45403 = ~w18568;
	assign w8502 = w45403 ^ w49450;
	assign w18459 = w18483 ^ w18460;
	assign w49442 = w18458 ^ w18459;
	assign w8243 = w49442 ^ w49446;
	assign w8521 = w8242 ^ w8243;
	assign w45626 = ~w27948;
	assign w45627 = ~w27949;
	assign w45628 = ~w27950;
	assign w45633 = ~w27947;
	assign w45710 = ~w31031;
	assign w45711 = ~w31032;
	assign w8203 = w8205 ^ w45711;
	assign w45716 = ~w31029;
	assign w8359 = w45716 ^ w45398;
	assign w45717 = ~w31030;
	assign w8467 = w45399 ^ w45717;
	assign w45920 = ~w7494;
	assign w7326 = w45920 ^ w45445;
	assign w48919 = w7326 ^ w7327;
	assign w7413 = w45920 ^ w49053;
	assign w47373 = w48919 ^ w1571;
	assign w19368 = w47376 ^ w47373;
	assign w19364 = w19368 ^ w19296;
	assign w19360 = w19279 ^ w19368;
	assign w19280 = w47375 ^ w47373;
	assign w19355 = w19280 ^ w19370;
	assign w19242 = w19282 ^ w19280;
	assign w19363 = w19280 ^ w19286;
	assign w19359 = w47380 ^ w19360;
	assign w19367 = w47373 ^ w47378;
	assign w19348 = w19363 & w19356;
	assign w19353 = w19360 & w19364;
	assign w19285 = w19353 ^ w19282;
	assign w19346 = w19370 & w19355;
	assign w19361 = w19296 ^ w19363;
	assign w7289 = w45920 ^ w49055;
	assign w19369 = w47373 ^ w47379;
	assign w19358 = w19279 ^ w19242;
	assign w19345 = w19367 & w19358;
	assign w7562 = w7289 ^ w7290;
	assign w48939 = w7562 ^ w7559;
	assign w47353 = w48939 ^ w1591;
	assign w31205 = w47355 ^ w47353;
	assign w31207 = w47354 ^ w31205;
	assign w31283 = w47350 ^ w31207;
	assign w31280 = w47351 ^ w31207;
	assign w31282 = w31212 ^ w31207;
	assign w31182 = w47353 ^ w47354;
	assign w31276 = w31295 & w31280;
	assign w31210 = w31276 ^ w31206;
	assign w31274 = w31289 & w31282;
	assign w19350 = w19369 & w19354;
	assign w44177 = w19345 ^ w19351;
	assign w44178 = w19345 ^ w19348;
	assign w19298 = w19346 ^ w44178;
	assign w19254 = w19349 ^ w19298;
	assign w19336 = w47379 ^ w19254;
	assign w19295 = w44177 ^ w19280;
	assign w48940 = w7412 ^ w7413;
	assign w47352 = w48940 ^ w1592;
	assign w31208 = w47352 ^ w47350;
	assign w31294 = w47352 ^ w47349;
	assign w31290 = w31294 ^ w31222;
	assign w31286 = w31205 ^ w31294;
	assign w31285 = w47356 ^ w31286;
	assign w31296 = w47354 ^ w47352;
	assign w31281 = w31206 ^ w31296;
	assign w31168 = w31208 ^ w31206;
	assign w31284 = w31205 ^ w31168;
	assign w31167 = w31208 ^ w47351;
	assign w31291 = w47356 ^ w31167;
	assign w31279 = w31286 & w31290;
	assign w31211 = w31279 ^ w31208;
	assign w31278 = w31287 & w31285;
	assign w31277 = w47356 & w31291;
	assign w31273 = w31294 & w31283;
	assign w31209 = w31273 ^ w31207;
	assign w31215 = w31211 ^ w31209;
	assign w31220 = w47349 ^ w31215;
	assign w31272 = w31296 & w31281;
	assign w31229 = w31272 ^ w31278;
	assign w31270 = w31229 ^ w31220;
	assign w31181 = w31272 ^ w31273;
	assign w31228 = w31181 ^ w31182;
	assign w31227 = w31228 ^ w31210;
	assign w31269 = w31275 ^ w31227;
	assign w31271 = w31293 & w31284;
	assign w31266 = w31270 & w31269;
	assign w44677 = w31271 ^ w31274;
	assign w31184 = w31210 ^ w44677;
	assign w31268 = w31184 ^ w31209;
	assign w31265 = w31266 ^ w31268;
	assign w31224 = w31272 ^ w44677;
	assign w31180 = w31275 ^ w31224;
	assign w31262 = w47355 ^ w31180;
	assign w44680 = w31271 ^ w31277;
	assign w31183 = w31215 ^ w44680;
	assign w31226 = w47351 ^ w31183;
	assign w31261 = w31266 ^ w31226;
	assign w31260 = w31261 & w31262;
	assign w31258 = w31266 ^ w31260;
	assign w31179 = w31260 ^ w31224;
	assign w31178 = w31260 ^ w31277;
	assign w31173 = w31178 ^ w31274;
	assign w31257 = w31268 & w31258;
	assign w31255 = w31257 ^ w31265;
	assign w44679 = w31257 ^ w31275;
	assign w31249 = w44679 ^ w31227;
	assign w31238 = w31249 & w31290;
	assign w31247 = w31249 & w31286;
	assign w31216 = w47355 ^ w44679;
	assign w31256 = w31216 ^ w31179;
	assign w31246 = w31256 & w31285;
	assign w31237 = w31256 & w31287;
	assign w31259 = w31260 ^ w31268;
	assign w31245 = w31259 & w47356;
	assign w31236 = w31259 & w31291;
	assign w31221 = w44680 ^ w31206;
	assign w31267 = w31229 ^ w31221;
	assign w31264 = w31267 & w31265;
	assign w31263 = w31264 ^ w31226;
	assign w31175 = w31264 ^ w31276;
	assign w31171 = w31175 ^ w31211;
	assign w31174 = w47349 ^ w31171;
	assign w31251 = w31173 ^ w31174;
	assign w31172 = w31264 ^ w31220;
	assign w31170 = w47351 ^ w31171;
	assign w31254 = w31263 & w31255;
	assign w31219 = w31254 ^ w31229;
	assign w31253 = w31219 ^ w31221;
	assign w31177 = w31254 ^ w31278;
	assign w31169 = w31216 ^ w31177;
	assign w31176 = w31206 ^ w31169;
	assign w31252 = w31173 ^ w31176;
	assign w31250 = w31219 ^ w31172;
	assign w31248 = w31169 ^ w31170;
	assign w31244 = w31250 & w31280;
	assign w31243 = w31253 & w31292;
	assign w31242 = w31263 & w31282;
	assign w31186 = w31242 ^ w31243;
	assign w31241 = w31251 & w31283;
	assign w31240 = w31248 & w31281;
	assign w31201 = w31240 ^ w31243;
	assign w31198 = ~w31201;
	assign w31197 = w31240 ^ w31241;
	assign w31239 = w31252 & w31284;
	assign w31235 = w31250 & w31295;
	assign w31217 = w31235 ^ w31239;
	assign w31202 = w31244 ^ w31235;
	assign w31195 = ~w31217;
	assign w31234 = w31253 & w31288;
	assign w31204 = w31242 ^ w31234;
	assign w31233 = w31263 & w31289;
	assign w31194 = w31195 ^ w31233;
	assign w31232 = w31251 & w31294;
	assign w31231 = w31248 & w31296;
	assign w31230 = w31252 & w31293;
	assign w31196 = w31241 ^ w31230;
	assign w31192 = ~w31196;
	assign w44678 = w31231 ^ w31232;
	assign w31213 = w31237 ^ w44678;
	assign w31214 = w31238 ^ w31213;
	assign w31218 = w31246 ^ w31214;
	assign w31187 = w31245 ^ w31218;
	assign w49257 = w31186 ^ w31187;
	assign w7724 = w49257 ^ w49247;
	assign w8028 = w49253 ^ w49257;
	assign w49124 = w8043 ^ w8028;
	assign w47241 = w49124 ^ w1703;
	assign w7908 = w7909 ^ w49257;
	assign w49132 = w7907 ^ w7908;
	assign w47233 = w49132 ^ w1711;
	assign w7893 = w8029 ^ w8028;
	assign w7891 = ~w7893;
	assign w31223 = w31247 ^ w31218;
	assign w31298 = w31223 ^ w31197;
	assign w7806 = w31298 ^ w49250;
	assign w49259 = ~w31298;
	assign w7900 = w8024 ^ w31298;
	assign w49135 = w7900 ^ w7901;
	assign w47230 = w49135 ^ w1714;
	assign w8018 = w45408 ^ w49259;
	assign w7825 = w8018 ^ w45641;
	assign w7916 = w8026 ^ w8018;
	assign w49127 = w45634 ^ w7916;
	assign w47238 = w49127 ^ w1706;
	assign w7887 = w8018 ^ w7974;
	assign w49144 = w49255 ^ w7887;
	assign w47221 = w49144 ^ w1723;
	assign w31200 = w31204 ^ w44678;
	assign w31199 = w31195 ^ w31200;
	assign w31299 = w31198 ^ w31199;
	assign w44681 = w31243 ^ w31244;
	assign w49258 = w44681 ^ w31223;
	assign w7843 = w49258 ^ w13073;
	assign w8025 = w49254 ^ w49258;
	assign w7890 = w8026 ^ w8025;
	assign w7918 = w7920 ^ w8025;
	assign w49142 = w45407 ^ w7890;
	assign w47223 = w49142 ^ w1721;
	assign w24640 = w47223 ^ w47221;
	assign w7760 = w7975 ^ w49258;
	assign w8045 = w7760 ^ w7761;
	assign w49133 = w8045 ^ w8029;
	assign w47232 = w49133 ^ w1712;
	assign w8104 = w47232 ^ w47230;
	assign w31225 = w31240 ^ w44681;
	assign w31191 = w31236 ^ w31225;
	assign w31188 = ~w31191;
	assign w31185 = w31241 ^ w31225;
	assign w49260 = w31214 ^ w31185;
	assign w7981 = w49244 ^ w49260;
	assign w7723 = w7981 ^ w49242;
	assign w8060 = w7723 ^ w7724;
	assign w7877 = ~w7981;
	assign w7876 = w7877 ^ w49246;
	assign w7973 = w49255 ^ w49260;
	assign w7897 = w8014 ^ w7973;
	assign w49117 = w8060 ^ w8025;
	assign w47248 = w49117 ^ w1696;
	assign w7966 = w8014 ^ w7981;
	assign w49137 = w45636 ^ w7897;
	assign w47228 = w49137 ^ w1716;
	assign w7915 = w8024 ^ w7973;
	assign w49128 = w49244 ^ w7915;
	assign w47237 = w49128 ^ w1707;
	assign w44682 = w31245 ^ w31247;
	assign w31203 = w44682 ^ w31200;
	assign w31300 = w31202 ^ w31203;
	assign w31190 = w31194 ^ w44682;
	assign w31193 = w31232 ^ w31190;
	assign w31297 = w31192 ^ w31193;
	assign w31189 = w31213 ^ w31190;
	assign w49256 = w31188 ^ w31189;
	assign w8016 = w49241 ^ w49256;
	assign w7878 = ~w8016;
	assign w7875 = w8028 ^ w7878;
	assign w49116 = w7875 ^ w7876;
	assign w47249 = w49116 ^ w1695;
	assign w7947 = w7878 ^ w45260;
	assign w49123 = w7947 ^ w7948;
	assign w47242 = w49123 ^ w1702;
	assign w12935 = w47237 ^ w47242;
	assign w12824 = w47241 ^ w47242;
	assign w7910 = w8016 ^ w8015;
	assign w49131 = w49245 ^ w7910;
	assign w47234 = w49131 ^ w1710;
	assign w8192 = w47234 ^ w47232;
	assign w8078 = w47233 ^ w47234;
	assign w19284 = w19350 ^ w19280;
	assign w19258 = w19284 ^ w44178;
	assign w19352 = w19361 & w19359;
	assign w19303 = w19346 ^ w19352;
	assign w19341 = w19303 ^ w19295;
	assign w45718 = ~w31299;
	assign w8036 = w45635 ^ w45718;
	assign w7889 = w8036 ^ w8013;
	assign w7912 = w8036 ^ w8014;
	assign w7906 = w7877 ^ w45718;
	assign w7895 = w45718 ^ w18703;
	assign w49115 = w49256 ^ w7889;
	assign w47250 = w49115 ^ w1694;
	assign w24864 = w47250 ^ w47248;
	assign w24750 = w47249 ^ w47250;
	assign w49139 = w7894 ^ w7895;
	assign w47226 = w49139 ^ w1718;
	assign w24727 = w47221 ^ w47226;
	assign w7911 = w7912 ^ w7913;
	assign w49130 = ~w7911;
	assign w47235 = w49130 ^ w1709;
	assign w8118 = w47235 ^ w47234;
	assign w8101 = w47235 ^ w47233;
	assign w8103 = w47234 ^ w8101;
	assign w8179 = w47230 ^ w8103;
	assign w45719 = ~w31300;
	assign w7766 = w7973 ^ w45719;
	assign w8042 = w7766 ^ w7767;
	assign w49138 = w8042 ^ w8015;
	assign w47227 = w49138 ^ w1717;
	assign w24656 = w47227 ^ w47226;
	assign w24729 = w47221 ^ w47227;
	assign w8037 = w45636 ^ w45719;
	assign w7789 = w8037 ^ w7974;
	assign w49121 = w45409 ^ w7789;
	assign w47244 = w49121 ^ w1700;
	assign w12854 = w47244 ^ w47238;
	assign w7914 = w8037 ^ w7975;
	assign w7905 = w8037 ^ w8015;
	assign w7904 = w7905 ^ w7906;
	assign w49114 = ~w7904;
	assign w47251 = w49114 ^ w1693;
	assign w24773 = w47251 ^ w47249;
	assign w24775 = w47250 ^ w24773;
	assign w24790 = w47251 ^ w47250;
	assign w49113 = w45719 ^ w7966;
	assign w47252 = w49113 ^ w1692;
	assign w49129 = w45261 ^ w7914;
	assign w47236 = w49129 ^ w1708;
	assign w8108 = w47236 ^ w47230;
	assign w8178 = w8108 ^ w8103;
	assign w45725 = ~w31297;
	assign w7902 = w8026 ^ w45725;
	assign w8021 = w45407 ^ w45725;
	assign w7888 = w8024 ^ w8021;
	assign w49134 = w7902 ^ w7903;
	assign w47231 = w49134 ^ w1713;
	assign w8188 = w47231 ^ w8108;
	assign w8176 = w47231 ^ w8103;
	assign w8184 = w47235 ^ w8188;
	assign w8171 = w8188 & w8184;
	assign w49143 = w45408 ^ w7888;
	assign w47222 = w49143 ^ w1722;
	assign w24646 = w47228 ^ w47222;
	assign w24723 = w24640 ^ w24646;
	assign w24721 = w24656 ^ w24723;
	assign w24726 = w47223 ^ w24646;
	assign w24722 = w47227 ^ w24726;
	assign w24709 = w24726 & w24722;
	assign w7826 = w45725 ^ w13074;
	assign w7824 = w7825 ^ w7826;
	assign w49119 = ~w7824;
	assign w47246 = w49119 ^ w1698;
	assign w24851 = w47246 ^ w24775;
	assign w24776 = w47248 ^ w47246;
	assign w24780 = w47252 ^ w47246;
	assign w24850 = w24780 ^ w24775;
	assign w7844 = w8021 ^ w49243;
	assign w7842 = ~w7844;
	assign w49118 = w7842 ^ w7843;
	assign w47247 = w49118 ^ w1697;
	assign w24848 = w47247 ^ w24775;
	assign w24860 = w47247 ^ w24780;
	assign w24856 = w47251 ^ w24860;
	assign w24735 = w24776 ^ w47247;
	assign w24859 = w47252 ^ w24735;
	assign w24845 = w47252 & w24859;
	assign w24843 = w24860 & w24856;
	assign w7917 = w8029 ^ w8021;
	assign w49126 = w45641 ^ w7917;
	assign w47239 = w49126 ^ w1705;
	assign w12934 = w47239 ^ w12854;
	assign w12848 = w47239 ^ w47237;
	assign w8063 = w8104 ^ w47231;
	assign w8187 = w47236 ^ w8063;
	assign w8173 = w47236 & w8187;
	assign w12931 = w12848 ^ w12854;
	assign w19347 = w19368 & w19357;
	assign w19255 = w19346 ^ w19347;
	assign w19302 = w19255 ^ w19256;
	assign w19301 = w19302 ^ w19284;
	assign w19343 = w19349 ^ w19301;
	assign w19283 = w19347 ^ w19281;
	assign w19342 = w19258 ^ w19283;
	assign w19289 = w19285 ^ w19283;
	assign w19257 = w19289 ^ w44177;
	assign w19300 = w47375 ^ w19257;
	assign w19294 = w47373 ^ w19289;
	assign w19344 = w19303 ^ w19294;
	assign w19340 = w19344 & w19343;
	assign w19335 = w19340 ^ w19300;
	assign w19334 = w19335 & w19336;
	assign w19253 = w19334 ^ w19298;
	assign w19333 = w19334 ^ w19342;
	assign w19310 = w19333 & w19365;
	assign w19319 = w19333 & w47380;
	assign w19332 = w19340 ^ w19334;
	assign w19331 = w19342 & w19332;
	assign w19339 = w19340 ^ w19342;
	assign w19338 = w19341 & w19339;
	assign w19249 = w19338 ^ w19350;
	assign w19329 = w19331 ^ w19339;
	assign w19337 = w19338 ^ w19300;
	assign w19328 = w19337 & w19329;
	assign w19251 = w19328 ^ w19352;
	assign w19293 = w19328 ^ w19303;
	assign w19327 = w19293 ^ w19295;
	assign w19308 = w19327 & w19362;
	assign w19317 = w19327 & w19366;
	assign w19252 = w19334 ^ w19351;
	assign w19247 = w19252 ^ w19348;
	assign w19245 = w19249 ^ w19285;
	assign w19248 = w47373 ^ w19245;
	assign w19325 = w19247 ^ w19248;
	assign w19246 = w19338 ^ w19294;
	assign w19324 = w19293 ^ w19246;
	assign w19309 = w19324 & w19369;
	assign w19318 = w19324 & w19354;
	assign w19276 = w19318 ^ w19309;
	assign w19316 = w19337 & w19356;
	assign w19278 = w19316 ^ w19308;
	assign w19315 = w19325 & w19357;
	assign w19307 = w19337 & w19363;
	assign w19306 = w19325 & w19368;
	assign w19244 = w47375 ^ w19245;
	assign w44179 = w19317 ^ w19318;
	assign w44181 = w19331 ^ w19349;
	assign w19323 = w44181 ^ w19301;
	assign w19321 = w19323 & w19360;
	assign w44180 = w19319 ^ w19321;
	assign w19312 = w19323 & w19364;
	assign w19290 = w47379 ^ w44181;
	assign w19243 = w19290 ^ w19251;
	assign w19330 = w19290 ^ w19253;
	assign w19311 = w19330 & w19361;
	assign w19320 = w19330 & w19359;
	assign w19250 = w19280 ^ w19243;
	assign w19326 = w19247 ^ w19250;
	assign w19304 = w19326 & w19367;
	assign w19270 = w19315 ^ w19304;
	assign w19313 = w19326 & w19358;
	assign w19266 = ~w19270;
	assign w19322 = w19243 ^ w19244;
	assign w19305 = w19322 & w19370;
	assign w19314 = w19322 & w19355;
	assign w19275 = w19314 ^ w19317;
	assign w19272 = ~w19275;
	assign w19299 = w19314 ^ w44179;
	assign w19259 = w19315 ^ w19299;
	assign w19265 = w19310 ^ w19299;
	assign w19271 = w19314 ^ w19315;
	assign w19262 = ~w19265;
	assign w43552 = w19305 ^ w19306;
	assign w19274 = w19278 ^ w43552;
	assign w19277 = w44180 ^ w19274;
	assign w19374 = w19276 ^ w19277;
	assign w19287 = w19311 ^ w43552;
	assign w19288 = w19312 ^ w19287;
	assign w49301 = w19288 ^ w19259;
	assign w19292 = w19320 ^ w19288;
	assign w19297 = w19321 ^ w19292;
	assign w49299 = w44179 ^ w19297;
	assign w19261 = w19319 ^ w19292;
	assign w7979 = w49301 ^ w49313;
	assign w7778 = w8017 ^ w7979;
	assign w49209 = w45259 ^ w7778;
	assign w47156 = w49209 ^ w1596;
	assign w7968 = w49301 ^ w49305;
	assign w7965 = w7979 ^ w49304;
	assign w8033 = w49299 ^ w49304;
	assign w49237 = w8039 ^ w8033;
	assign w47128 = w49237 ^ w1624;
	assign w7938 = w8033 ^ w7987;
	assign w7773 = ~w49299;
	assign w7772 = w49303 ^ w7773;
	assign w7962 = w49312 ^ w7773;
	assign w49214 = w7961 ^ w7962;
	assign w7957 = w8017 ^ w7968;
	assign w49229 = w7938 ^ w7939;
	assign w7933 = w7968 ^ w49313;
	assign w49232 = w7933 ^ w7934;
	assign w47133 = w49232 ^ w1619;
	assign w47151 = w49214 ^ w1601;
	assign w47136 = w49229 ^ w1616;
	assign w19372 = w19297 ^ w19271;
	assign w49300 = ~w19372;
	assign w8032 = w49300 ^ w45265;
	assign w7922 = w8032 ^ w45200;
	assign w7943 = w8032 ^ w7967;
	assign w7959 = w49305 ^ w19372;
	assign w49224 = w49301 ^ w7943;
	assign w7935 = w8032 ^ w7992;
	assign w49231 = w45197 ^ w7935;
	assign w47141 = w49224 ^ w1611;
	assign w47134 = w49231 ^ w1618;
	assign w18076 = w47136 ^ w47134;
	assign w49239 = w7922 ^ w7923;
	assign w47126 = w49239 ^ w1626;
	assign w24508 = w47128 ^ w47126;
	assign w7921 = w7990 ^ w7968;
	assign w49240 = w49309 ^ w7921;
	assign w47125 = w49240 ^ w1627;
	assign w24594 = w47128 ^ w47125;
	assign w19291 = w19309 ^ w19313;
	assign w19269 = ~w19291;
	assign w19273 = w19269 ^ w19274;
	assign w19373 = w19272 ^ w19273;
	assign w19268 = w19269 ^ w19307;
	assign w19264 = w19268 ^ w44180;
	assign w19267 = w19306 ^ w19264;
	assign w19371 = w19266 ^ w19267;
	assign w19263 = w19287 ^ w19264;
	assign w18162 = w47136 ^ w47133;
	assign w49297 = w19262 ^ w19263;
	assign w7735 = w7979 ^ w49297;
	assign w8055 = w7735 ^ w7736;
	assign w49212 = w8055 ^ w7987;
	assign w47153 = w49212 ^ w1599;
	assign w8007 = w49297 ^ w49302;
	assign w7928 = w8007 ^ w7997;
	assign w7940 = w8007 ^ w49310;
	assign w49227 = w7940 ^ w7941;
	assign w47138 = w49227 ^ w1614;
	assign w18164 = w47138 ^ w47136;
	assign w18161 = w47133 ^ w47138;
	assign w49235 = w49306 ^ w7928;
	assign w47130 = w49235 ^ w1622;
	assign w24596 = w47130 ^ w47128;
	assign w24593 = w47125 ^ w47130;
	assign w45422 = ~w19374;
	assign w7733 = w7979 ^ w45422;
	assign w8056 = w7733 ^ w7734;
	assign w49210 = w8056 ^ w7997;
	assign w8030 = w45422 ^ w45259;
	assign w7955 = w8030 ^ w7997;
	assign w7942 = w8030 ^ w7982;
	assign w49225 = w45199 ^ w7942;
	assign w47140 = w49225 ^ w1612;
	assign w18080 = w47140 ^ w47134;
	assign w7932 = w8030 ^ w7967;
	assign w49233 = w45632 ^ w7932;
	assign w47132 = w49233 ^ w1620;
	assign w24512 = w47132 ^ w47126;
	assign w47155 = w49210 ^ w1597;
	assign w27721 = w47155 ^ w47153;
	assign w49217 = w45422 ^ w7957;
	assign w47148 = w49217 ^ w1604;
	assign w45428 = ~w19371;
	assign w7946 = w19372 ^ w45428;
	assign w7944 = w7945 ^ w7946;
	assign w49223 = ~w7944;
	assign w49238 = w45428 ^ w7924;
	assign w47127 = w49238 ^ w1625;
	assign w24506 = w47127 ^ w47125;
	assign w24581 = w24506 ^ w24596;
	assign w24589 = w24506 ^ w24512;
	assign w24592 = w47127 ^ w24512;
	assign w24468 = w24508 ^ w24506;
	assign w24467 = w24508 ^ w47127;
	assign w24591 = w47132 ^ w24467;
	assign w24577 = w47132 & w24591;
	assign w24572 = w24596 & w24581;
	assign w47142 = w49223 ^ w1610;
	assign w12586 = w47148 ^ w47142;
	assign w8002 = w45428 ^ w45200;
	assign w7936 = w8002 ^ w49308;
	assign w49230 = w7936 ^ w7937;
	assign w7949 = w8033 ^ w8002;
	assign w49222 = w45637 ^ w7949;
	assign w7960 = w8002 ^ w7990;
	assign w47143 = w49222 ^ w1609;
	assign w12666 = w47143 ^ w12586;
	assign w47135 = w49230 ^ w1617;
	assign w18074 = w47135 ^ w47133;
	assign w18149 = w18074 ^ w18164;
	assign w18160 = w47135 ^ w18080;
	assign w18157 = w18074 ^ w18080;
	assign w18036 = w18076 ^ w18074;
	assign w18140 = w18164 & w18149;
	assign w18035 = w18076 ^ w47135;
	assign w18159 = w47140 ^ w18035;
	assign w18145 = w47140 & w18159;
	assign w12580 = w47143 ^ w47141;
	assign w12663 = w12580 ^ w12586;
	assign w49215 = w45265 ^ w7960;
	assign w47150 = w49215 ^ w1602;
	assign w27728 = w47156 ^ w47150;
	assign w27808 = w47151 ^ w27728;
	assign w27804 = w47155 ^ w27808;
	assign w27791 = w27808 & w27804;
	assign w45429 = ~w19373;
	assign w7776 = w7985 ^ w45429;
	assign w49211 = w7776 ^ w7777;
	assign w8022 = w45429 ^ w45258;
	assign w49226 = w8062 ^ w8022;
	assign w7931 = ~w8022;
	assign w7929 = w7931 ^ w8017;
	assign w7953 = w8022 ^ w7985;
	assign w49219 = w49297 ^ w7953;
	assign w47146 = w49219 ^ w1606;
	assign w12667 = w47141 ^ w47146;
	assign w47139 = w49226 ^ w1613;
	assign w18090 = w47139 ^ w47138;
	assign w18155 = w18090 ^ w18157;
	assign w18156 = w47139 ^ w18160;
	assign w18158 = w18162 ^ w18090;
	assign w18143 = w18160 & w18156;
	assign w18163 = w47133 ^ w47139;
	assign w47154 = w49211 ^ w1598;
	assign w27723 = w47154 ^ w27721;
	assign w27799 = w47150 ^ w27723;
	assign w27796 = w47151 ^ w27723;
	assign w27798 = w27728 ^ w27723;
	assign w27738 = w47155 ^ w47154;
	assign w27698 = w47153 ^ w47154;
	assign w19260 = w19316 ^ w19317;
	assign w49298 = w19260 ^ w19261;
	assign w7993 = w49298 ^ w49311;
	assign w49228 = w8061 ^ w7993;
	assign w7952 = w8007 ^ w7993;
	assign w7950 = ~w7952;
	assign w7964 = w7993 ^ w7984;
	assign w49213 = w7964 ^ w7965;
	assign w47152 = w49213 ^ w1600;
	assign w27724 = w47152 ^ w47150;
	assign w27812 = w47154 ^ w47152;
	assign w27683 = w27724 ^ w47151;
	assign w27807 = w47156 ^ w27683;
	assign w27793 = w47156 & w27807;
	assign w47137 = w49228 ^ w1615;
	assign w18050 = w47137 ^ w47138;
	assign w18073 = w47139 ^ w47137;
	assign w18154 = w18073 ^ w18162;
	assign w18153 = w47140 ^ w18154;
	assign w18075 = w47138 ^ w18073;
	assign w18148 = w47135 ^ w18075;
	assign w18151 = w47134 ^ w18075;
	assign w18150 = w18080 ^ w18075;
	assign w18152 = w18073 ^ w18036;
	assign w18146 = w18155 & w18153;
	assign w18144 = w18163 & w18148;
	assign w18078 = w18144 ^ w18074;
	assign w18147 = w18154 & w18158;
	assign w18079 = w18147 ^ w18076;
	assign w18142 = w18157 & w18150;
	assign w18141 = w18162 & w18151;
	assign w18049 = w18140 ^ w18141;
	assign w18096 = w18049 ^ w18050;
	assign w18095 = w18096 ^ w18078;
	assign w18137 = w18143 ^ w18095;
	assign w18077 = w18141 ^ w18075;
	assign w18083 = w18079 ^ w18077;
	assign w18088 = w47133 ^ w18083;
	assign w18139 = w18161 & w18152;
	assign w44126 = w18139 ^ w18145;
	assign w18089 = w44126 ^ w18074;
	assign w18051 = w18083 ^ w44126;
	assign w18094 = w47135 ^ w18051;
	assign w44127 = w18139 ^ w18142;
	assign w18092 = w18140 ^ w44127;
	assign w18048 = w18143 ^ w18092;
	assign w18130 = w47139 ^ w18048;
	assign w18052 = w18078 ^ w44127;
	assign w18136 = w18052 ^ w18077;
	assign w18097 = w18140 ^ w18146;
	assign w18138 = w18097 ^ w18088;
	assign w18134 = w18138 & w18137;
	assign w18129 = w18134 ^ w18094;
	assign w18128 = w18129 & w18130;
	assign w18126 = w18134 ^ w18128;
	assign w18047 = w18128 ^ w18092;
	assign w18127 = w18128 ^ w18136;
	assign w18113 = w18127 & w47140;
	assign w18104 = w18127 & w18159;
	assign w18125 = w18136 & w18126;
	assign w44130 = w18125 ^ w18143;
	assign w18084 = w47139 ^ w44130;
	assign w18124 = w18084 ^ w18047;
	assign w18114 = w18124 & w18153;
	assign w18105 = w18124 & w18155;
	assign w18117 = w44130 ^ w18095;
	assign w18106 = w18117 & w18158;
	assign w18115 = w18117 & w18154;
	assign w44129 = w18113 ^ w18115;
	assign w18046 = w18128 ^ w18145;
	assign w18041 = w18046 ^ w18142;
	assign w18135 = w18097 ^ w18089;
	assign w18133 = w18134 ^ w18136;
	assign w18123 = w18125 ^ w18133;
	assign w18132 = w18135 & w18133;
	assign w18131 = w18132 ^ w18094;
	assign w18110 = w18131 & w18150;
	assign w18043 = w18132 ^ w18144;
	assign w18040 = w18132 ^ w18088;
	assign w18039 = w18043 ^ w18079;
	assign w18042 = w47133 ^ w18039;
	assign w18119 = w18041 ^ w18042;
	assign w18100 = w18119 & w18162;
	assign w18109 = w18119 & w18151;
	assign w18038 = w47135 ^ w18039;
	assign w18101 = w18131 & w18157;
	assign w18122 = w18131 & w18123;
	assign w18087 = w18122 ^ w18097;
	assign w18118 = w18087 ^ w18040;
	assign w18103 = w18118 & w18163;
	assign w18121 = w18087 ^ w18089;
	assign w18045 = w18122 ^ w18146;
	assign w18037 = w18084 ^ w18045;
	assign w18044 = w18074 ^ w18037;
	assign w18102 = w18121 & w18156;
	assign w18072 = w18110 ^ w18102;
	assign w18120 = w18041 ^ w18044;
	assign w18111 = w18121 & w18160;
	assign w18054 = w18110 ^ w18111;
	assign w18116 = w18037 ^ w18038;
	assign w18099 = w18116 & w18164;
	assign w18107 = w18120 & w18152;
	assign w18108 = w18116 & w18149;
	assign w18069 = w18108 ^ w18111;
	assign w18066 = ~w18069;
	assign w18065 = w18108 ^ w18109;
	assign w18098 = w18120 & w18161;
	assign w18064 = w18109 ^ w18098;
	assign w18060 = ~w18064;
	assign w43549 = w18099 ^ w18100;
	assign w18081 = w18105 ^ w43549;
	assign w18082 = w18106 ^ w18081;
	assign w18086 = w18114 ^ w18082;
	assign w18055 = w18113 ^ w18086;
	assign w49454 = w18054 ^ w18055;
	assign w8239 = w49454 ^ w49447;
	assign w18091 = w18115 ^ w18086;
	assign w18068 = w18072 ^ w43549;
	assign w18071 = w44129 ^ w18068;
	assign w18112 = w18118 & w18148;
	assign w18070 = w18112 ^ w18103;
	assign w18168 = w18070 ^ w18071;
	assign w44128 = w18111 ^ w18112;
	assign w18093 = w18108 ^ w44128;
	assign w18059 = w18104 ^ w18093;
	assign w18056 = ~w18059;
	assign w18053 = w18109 ^ w18093;
	assign w49456 = w18082 ^ w18053;
	assign w8453 = w49451 ^ w49456;
	assign w8387 = ~w8453;
	assign w8391 = w8387 ^ w45779;
	assign w49455 = w44128 ^ w18091;
	assign w8381 = w49455 ^ w49448;
	assign w18085 = w18103 ^ w18107;
	assign w18063 = ~w18085;
	assign w18062 = w18063 ^ w18101;
	assign w18058 = w18062 ^ w44129;
	assign w18061 = w18100 ^ w18058;
	assign w18165 = w18060 ^ w18061;
	assign w18057 = w18081 ^ w18058;
	assign w49453 = w18056 ^ w18057;
	assign w8491 = w49446 ^ w49453;
	assign w8374 = ~w8491;
	assign w8385 = w8516 ^ w8374;
	assign w8248 = ~w49453;
	assign w8247 = w49454 ^ w8248;
	assign w8426 = w45404 ^ w8248;
	assign w8372 = w8374 ^ w49442;
	assign w18067 = w18063 ^ w18068;
	assign w18167 = w18066 ^ w18067;
	assign w49452 = ~w18167;
	assign w8493 = w45779 ^ w49452;
	assign w8241 = w18167 ^ w45405;
	assign w18166 = w18091 ^ w18065;
	assign w45390 = ~w18165;
	assign w8379 = w45390 ^ w33709;
	assign w45391 = ~w18166;
	assign w8377 = w45391 ^ w33710;
	assign w45392 = ~w18168;
	assign w8492 = w45780 ^ w45392;
	assign w8245 = w45404 ^ w45392;
	assign w45921 = ~w7968;
	assign w7771 = w45921 ^ w49298;
	assign w8040 = w7771 ^ w7772;
	assign w49221 = w8040 ^ w7984;
	assign w7956 = w45921 ^ w45429;
	assign w7951 = w45921 ^ w49307;
	assign w49220 = w7950 ^ w7951;
	assign w47145 = w49220 ^ w1607;
	assign w12556 = w47145 ^ w47146;
	assign w7954 = w7955 ^ w7956;
	assign w49218 = ~w7954;
	assign w47144 = w49221 ^ w1608;
	assign w12582 = w47144 ^ w47142;
	assign w12541 = w12582 ^ w47143;
	assign w12665 = w47148 ^ w12541;
	assign w12542 = w12582 ^ w12580;
	assign w12651 = w47148 & w12665;
	assign w12668 = w47144 ^ w47141;
	assign w12670 = w47146 ^ w47144;
	assign w47147 = w49218 ^ w1605;
	assign w12579 = w47147 ^ w47145;
	assign w12669 = w47141 ^ w47147;
	assign w12658 = w12579 ^ w12542;
	assign w12645 = w12667 & w12658;
	assign w12660 = w12579 ^ w12668;
	assign w12596 = w47147 ^ w47146;
	assign w12664 = w12668 ^ w12596;
	assign w12661 = w12596 ^ w12663;
	assign w12662 = w47147 ^ w12666;
	assign w12649 = w12666 & w12662;
	assign w12659 = w47148 ^ w12660;
	assign w12652 = w12661 & w12659;
	assign w12655 = w12580 ^ w12670;
	assign w12646 = w12670 & w12655;
	assign w12603 = w12646 ^ w12652;
	assign w43897 = w12645 ^ w12651;
	assign w12595 = w43897 ^ w12580;
	assign w12641 = w12603 ^ w12595;
	assign w12581 = w47146 ^ w12579;
	assign w12657 = w47142 ^ w12581;
	assign w12647 = w12668 & w12657;
	assign w12583 = w12647 ^ w12581;
	assign w12555 = w12646 ^ w12647;
	assign w12654 = w47143 ^ w12581;
	assign w12650 = w12669 & w12654;
	assign w12584 = w12650 ^ w12580;
	assign w12656 = w12586 ^ w12581;
	assign w12648 = w12663 & w12656;
	assign w12602 = w12555 ^ w12556;
	assign w12601 = w12602 ^ w12584;
	assign w12643 = w12649 ^ w12601;
	assign w12653 = w12660 & w12664;
	assign w12585 = w12653 ^ w12582;
	assign w12589 = w12585 ^ w12583;
	assign w12557 = w12589 ^ w43897;
	assign w12600 = w47143 ^ w12557;
	assign w12594 = w47141 ^ w12589;
	assign w12644 = w12603 ^ w12594;
	assign w12640 = w12644 & w12643;
	assign w12635 = w12640 ^ w12600;
	assign w43898 = w12645 ^ w12648;
	assign w12558 = w12584 ^ w43898;
	assign w12642 = w12558 ^ w12583;
	assign w12639 = w12640 ^ w12642;
	assign w12638 = w12641 & w12639;
	assign w12549 = w12638 ^ w12650;
	assign w12545 = w12549 ^ w12585;
	assign w12548 = w47141 ^ w12545;
	assign w12544 = w47143 ^ w12545;
	assign w12637 = w12638 ^ w12600;
	assign w12607 = w12637 & w12663;
	assign w12616 = w12637 & w12656;
	assign w12546 = w12638 ^ w12594;
	assign w12598 = w12646 ^ w43898;
	assign w12554 = w12649 ^ w12598;
	assign w12636 = w47147 ^ w12554;
	assign w12634 = w12635 & w12636;
	assign w12552 = w12634 ^ w12651;
	assign w12553 = w12634 ^ w12598;
	assign w12632 = w12640 ^ w12634;
	assign w12631 = w12642 & w12632;
	assign w12633 = w12634 ^ w12642;
	assign w12610 = w12633 & w12665;
	assign w12629 = w12631 ^ w12639;
	assign w12628 = w12637 & w12629;
	assign w12551 = w12628 ^ w12652;
	assign w12593 = w12628 ^ w12603;
	assign w12624 = w12593 ^ w12546;
	assign w12609 = w12624 & w12669;
	assign w12627 = w12593 ^ w12595;
	assign w12608 = w12627 & w12662;
	assign w12578 = w12616 ^ w12608;
	assign w12619 = w12633 & w47148;
	assign w12618 = w12624 & w12654;
	assign w12576 = w12618 ^ w12609;
	assign w12547 = w12552 ^ w12648;
	assign w12625 = w12547 ^ w12548;
	assign w12615 = w12625 & w12657;
	assign w12606 = w12625 & w12668;
	assign w43902 = w12631 ^ w12649;
	assign w12623 = w43902 ^ w12601;
	assign w12612 = w12623 & w12664;
	assign w12621 = w12623 & w12660;
	assign w43901 = w12619 ^ w12621;
	assign w12590 = w47147 ^ w43902;
	assign w12543 = w12590 ^ w12551;
	assign w12622 = w12543 ^ w12544;
	assign w12550 = w12580 ^ w12543;
	assign w12605 = w12622 & w12670;
	assign w12626 = w12547 ^ w12550;
	assign w12604 = w12626 & w12667;
	assign w12613 = w12626 & w12658;
	assign w12570 = w12615 ^ w12604;
	assign w12566 = ~w12570;
	assign w12591 = w12609 ^ w12613;
	assign w12569 = ~w12591;
	assign w12568 = w12569 ^ w12607;
	assign w12564 = w12568 ^ w43901;
	assign w12567 = w12606 ^ w12564;
	assign w12671 = w12566 ^ w12567;
	assign w43899 = w12605 ^ w12606;
	assign w12574 = w12578 ^ w43899;
	assign w12577 = w43901 ^ w12574;
	assign w12573 = w12569 ^ w12574;
	assign w12674 = w12576 ^ w12577;
	assign w12617 = w12627 & w12666;
	assign w12560 = w12616 ^ w12617;
	assign w43900 = w12617 ^ w12618;
	assign w12614 = w12622 & w12655;
	assign w12571 = w12614 ^ w12615;
	assign w12575 = w12614 ^ w12617;
	assign w12572 = ~w12575;
	assign w12599 = w12614 ^ w43900;
	assign w12559 = w12615 ^ w12599;
	assign w12673 = w12572 ^ w12573;
	assign w8204 = w12673 ^ w45401;
	assign w8537 = w8203 ^ w8204;
	assign w49466 = ~w12673;
	assign w8488 = w45400 ^ w49466;
	assign w12565 = w12610 ^ w12599;
	assign w12562 = ~w12565;
	assign w45251 = ~w12671;
	assign w8361 = w45251 ^ w49464;
	assign w8473 = w45398 ^ w45251;
	assign w8341 = w8473 ^ w8467;
	assign w8334 = w8473 ^ w45716;
	assign w8332 = ~w8334;
	assign w45253 = ~w12674;
	assign w8489 = w45401 ^ w45253;
	assign w12630 = w12590 ^ w12553;
	assign w12611 = w12630 & w12661;
	assign w12620 = w12630 & w12659;
	assign w12587 = w12611 ^ w43899;
	assign w12563 = w12587 ^ w12564;
	assign w49467 = w12562 ^ w12563;
	assign w8363 = w49467 ^ w45400;
	assign w8484 = w49462 ^ w49467;
	assign w8337 = ~w8484;
	assign w8335 = w8337 ^ w49475;
	assign w12588 = w12612 ^ w12587;
	assign w49470 = w12588 ^ w12559;
	assign w8449 = w49465 ^ w49470;
	assign w8312 = w8449 ^ w45717;
	assign w12592 = w12620 ^ w12588;
	assign w12561 = w12619 ^ w12592;
	assign w12597 = w12621 ^ w12592;
	assign w12672 = w12597 ^ w12571;
	assign w49468 = w12560 ^ w12561;
	assign w8208 = ~w49468;
	assign w8207 = w8208 ^ w49462;
	assign w8536 = w8206 ^ w8207;
	assign w8481 = w49463 ^ w49468;
	assign w8345 = ~w8481;
	assign w49469 = w43900 ^ w12597;
	assign w8210 = w49469 ^ w49463;
	assign w8535 = w8209 ^ w8210;
	assign w8477 = w49464 ^ w49469;
	assign w8319 = ~w8477;
	assign w45252 = ~w12672;
	assign w8331 = w45252 ^ w45251;
	assign w45922 = ~w7967;
	assign w7958 = w45922 ^ w45197;
	assign w7930 = w45922 ^ w45631;
	assign w49234 = w7929 ^ w7930;
	assign w7927 = w45922 ^ w49298;
	assign w49216 = w7958 ^ w7959;
	assign w47149 = w49216 ^ w1603;
	assign w27722 = w47151 ^ w47149;
	assign w27797 = w27722 ^ w27812;
	assign w27810 = w47152 ^ w47149;
	assign w27806 = w27810 ^ w27738;
	assign w27805 = w27722 ^ w27728;
	assign w27803 = w27738 ^ w27805;
	assign w27802 = w27721 ^ w27810;
	assign w27801 = w47156 ^ w27802;
	assign w27684 = w27724 ^ w27722;
	assign w27800 = w27721 ^ w27684;
	assign w27811 = w47149 ^ w47155;
	assign w27809 = w47149 ^ w47154;
	assign w27795 = w27802 & w27806;
	assign w27727 = w27795 ^ w27724;
	assign w27794 = w27803 & w27801;
	assign w27792 = w27811 & w27796;
	assign w27726 = w27792 ^ w27722;
	assign w27790 = w27805 & w27798;
	assign w27789 = w27810 & w27799;
	assign w27725 = w27789 ^ w27723;
	assign w27731 = w27727 ^ w27725;
	assign w27736 = w47149 ^ w27731;
	assign w27788 = w27812 & w27797;
	assign w27745 = w27788 ^ w27794;
	assign w27786 = w27745 ^ w27736;
	assign w27697 = w27788 ^ w27789;
	assign w27744 = w27697 ^ w27698;
	assign w27743 = w27744 ^ w27726;
	assign w27785 = w27791 ^ w27743;
	assign w27787 = w27809 & w27800;
	assign w27782 = w27786 & w27785;
	assign w7925 = w7926 ^ w7927;
	assign w49236 = ~w7925;
	assign w47129 = w49236 ^ w1623;
	assign w24482 = w47129 ^ w47130;
	assign w47131 = w49234 ^ w1621;
	assign w24505 = w47131 ^ w47129;
	assign w24507 = w47130 ^ w24505;
	assign w24583 = w47126 ^ w24507;
	assign w24580 = w47127 ^ w24507;
	assign w24582 = w24512 ^ w24507;
	assign w24588 = w47131 ^ w24592;
	assign w24586 = w24505 ^ w24594;
	assign w24585 = w47132 ^ w24586;
	assign w24522 = w47131 ^ w47130;
	assign w24587 = w24522 ^ w24589;
	assign w24590 = w24594 ^ w24522;
	assign w24584 = w24505 ^ w24468;
	assign w24595 = w47125 ^ w47131;
	assign w24579 = w24586 & w24590;
	assign w24511 = w24579 ^ w24508;
	assign w24578 = w24587 & w24585;
	assign w24529 = w24572 ^ w24578;
	assign w24576 = w24595 & w24580;
	assign w24510 = w24576 ^ w24506;
	assign w24575 = w24592 & w24588;
	assign w24574 = w24589 & w24582;
	assign w24573 = w24594 & w24583;
	assign w24509 = w24573 ^ w24507;
	assign w24515 = w24511 ^ w24509;
	assign w24520 = w47125 ^ w24515;
	assign w24570 = w24529 ^ w24520;
	assign w24481 = w24572 ^ w24573;
	assign w24528 = w24481 ^ w24482;
	assign w24527 = w24528 ^ w24510;
	assign w24569 = w24575 ^ w24527;
	assign w24571 = w24593 & w24584;
	assign w24566 = w24570 & w24569;
	assign w44396 = w24571 ^ w24577;
	assign w24483 = w24515 ^ w44396;
	assign w24526 = w47127 ^ w24483;
	assign w24561 = w24566 ^ w24526;
	assign w24521 = w44396 ^ w24506;
	assign w24567 = w24529 ^ w24521;
	assign w44397 = w24571 ^ w24574;
	assign w24524 = w24572 ^ w44397;
	assign w24480 = w24575 ^ w24524;
	assign w24562 = w47131 ^ w24480;
	assign w24560 = w24561 & w24562;
	assign w24558 = w24566 ^ w24560;
	assign w24479 = w24560 ^ w24524;
	assign w24478 = w24560 ^ w24577;
	assign w24473 = w24478 ^ w24574;
	assign w24484 = w24510 ^ w44397;
	assign w24568 = w24484 ^ w24509;
	assign w24559 = w24560 ^ w24568;
	assign w24565 = w24566 ^ w24568;
	assign w24564 = w24567 & w24565;
	assign w24563 = w24564 ^ w24526;
	assign w24475 = w24564 ^ w24576;
	assign w24471 = w24475 ^ w24511;
	assign w24474 = w47125 ^ w24471;
	assign w24551 = w24473 ^ w24474;
	assign w24472 = w24564 ^ w24520;
	assign w24470 = w47127 ^ w24471;
	assign w24557 = w24568 & w24558;
	assign w24555 = w24557 ^ w24565;
	assign w24554 = w24563 & w24555;
	assign w24519 = w24554 ^ w24529;
	assign w24553 = w24519 ^ w24521;
	assign w24477 = w24554 ^ w24578;
	assign w24550 = w24519 ^ w24472;
	assign w24545 = w24559 & w47132;
	assign w24544 = w24550 & w24580;
	assign w24543 = w24553 & w24592;
	assign w24542 = w24563 & w24582;
	assign w24486 = w24542 ^ w24543;
	assign w24541 = w24551 & w24583;
	assign w24536 = w24559 & w24591;
	assign w24535 = w24550 & w24595;
	assign w24502 = w24544 ^ w24535;
	assign w24534 = w24553 & w24588;
	assign w24504 = w24542 ^ w24534;
	assign w24533 = w24563 & w24589;
	assign w24532 = w24551 & w24594;
	assign w44399 = w24543 ^ w24544;
	assign w44401 = w24557 ^ w24575;
	assign w24549 = w44401 ^ w24527;
	assign w24538 = w24549 & w24590;
	assign w24547 = w24549 & w24586;
	assign w44400 = w24545 ^ w24547;
	assign w24516 = w47131 ^ w44401;
	assign w24556 = w24516 ^ w24479;
	assign w24469 = w24516 ^ w24477;
	assign w24476 = w24506 ^ w24469;
	assign w24552 = w24473 ^ w24476;
	assign w24548 = w24469 ^ w24470;
	assign w24546 = w24556 & w24585;
	assign w24540 = w24548 & w24581;
	assign w24525 = w24540 ^ w44399;
	assign w24501 = w24540 ^ w24543;
	assign w24498 = ~w24501;
	assign w24497 = w24540 ^ w24541;
	assign w24491 = w24536 ^ w24525;
	assign w24488 = ~w24491;
	assign w24485 = w24541 ^ w24525;
	assign w24539 = w24552 & w24584;
	assign w24517 = w24535 ^ w24539;
	assign w24495 = ~w24517;
	assign w24494 = w24495 ^ w24533;
	assign w24490 = w24494 ^ w44400;
	assign w24493 = w24532 ^ w24490;
	assign w24537 = w24556 & w24587;
	assign w24531 = w24548 & w24596;
	assign w24530 = w24552 & w24593;
	assign w24496 = w24541 ^ w24530;
	assign w24492 = ~w24496;
	assign w24597 = w24492 ^ w24493;
	assign w44398 = w24531 ^ w24532;
	assign w24513 = w24537 ^ w44398;
	assign w24514 = w24538 ^ w24513;
	assign w24518 = w24546 ^ w24514;
	assign w24523 = w24547 ^ w24518;
	assign w49513 = w44399 ^ w24523;
	assign w8462 = w49509 ^ w49513;
	assign w24598 = w24523 ^ w24497;
	assign w24489 = w24513 ^ w24490;
	assign w49511 = w24488 ^ w24489;
	assign w24487 = w24545 ^ w24518;
	assign w49512 = w24486 ^ w24487;
	assign w49514 = w24514 ^ w24485;
	assign w8445 = w49510 ^ w49514;
	assign w8214 = w49512 ^ w49511;
	assign w8252 = w8445 ^ w49512;
	assign w8517 = w8252 ^ w8253;
	assign w8463 = w49507 ^ w49511;
	assign w24500 = w24504 ^ w44398;
	assign w24503 = w44400 ^ w24500;
	assign w24600 = w24502 ^ w24503;
	assign w24499 = w24495 ^ w24500;
	assign w24599 = w24498 ^ w24499;
	assign w44528 = w27787 ^ w27793;
	assign w27699 = w27731 ^ w44528;
	assign w27742 = w47151 ^ w27699;
	assign w27777 = w27782 ^ w27742;
	assign w27737 = w44528 ^ w27722;
	assign w27783 = w27745 ^ w27737;
	assign w44529 = w27787 ^ w27790;
	assign w27740 = w27788 ^ w44529;
	assign w27696 = w27791 ^ w27740;
	assign w27778 = w47155 ^ w27696;
	assign w27776 = w27777 & w27778;
	assign w27774 = w27782 ^ w27776;
	assign w27695 = w27776 ^ w27740;
	assign w27694 = w27776 ^ w27793;
	assign w27689 = w27694 ^ w27790;
	assign w27700 = w27726 ^ w44529;
	assign w27784 = w27700 ^ w27725;
	assign w27775 = w27776 ^ w27784;
	assign w27781 = w27782 ^ w27784;
	assign w27780 = w27783 & w27781;
	assign w27779 = w27780 ^ w27742;
	assign w27691 = w27780 ^ w27792;
	assign w27687 = w27691 ^ w27727;
	assign w27690 = w47149 ^ w27687;
	assign w27767 = w27689 ^ w27690;
	assign w27688 = w27780 ^ w27736;
	assign w27686 = w47151 ^ w27687;
	assign w27773 = w27784 & w27774;
	assign w27771 = w27773 ^ w27781;
	assign w27770 = w27779 & w27771;
	assign w27735 = w27770 ^ w27745;
	assign w27769 = w27735 ^ w27737;
	assign w27693 = w27770 ^ w27794;
	assign w27766 = w27735 ^ w27688;
	assign w27761 = w27775 & w47156;
	assign w27760 = w27766 & w27796;
	assign w27759 = w27769 & w27808;
	assign w27758 = w27779 & w27798;
	assign w27702 = w27758 ^ w27759;
	assign w27757 = w27767 & w27799;
	assign w27752 = w27775 & w27807;
	assign w27751 = w27766 & w27811;
	assign w27718 = w27760 ^ w27751;
	assign w27750 = w27769 & w27804;
	assign w27720 = w27758 ^ w27750;
	assign w27749 = w27779 & w27805;
	assign w27748 = w27767 & w27810;
	assign w44531 = w27759 ^ w27760;
	assign w44533 = w27773 ^ w27791;
	assign w27765 = w44533 ^ w27743;
	assign w27763 = w27765 & w27802;
	assign w44532 = w27761 ^ w27763;
	assign w27754 = w27765 & w27806;
	assign w27732 = w47155 ^ w44533;
	assign w27772 = w27732 ^ w27695;
	assign w27685 = w27732 ^ w27693;
	assign w27692 = w27722 ^ w27685;
	assign w27768 = w27689 ^ w27692;
	assign w27764 = w27685 ^ w27686;
	assign w27762 = w27772 & w27801;
	assign w27756 = w27764 & w27797;
	assign w27741 = w27756 ^ w44531;
	assign w27717 = w27756 ^ w27759;
	assign w27714 = ~w27717;
	assign w27713 = w27756 ^ w27757;
	assign w27707 = w27752 ^ w27741;
	assign w27704 = ~w27707;
	assign w27701 = w27757 ^ w27741;
	assign w27755 = w27768 & w27800;
	assign w27733 = w27751 ^ w27755;
	assign w27711 = ~w27733;
	assign w27710 = w27711 ^ w27749;
	assign w27706 = w27710 ^ w44532;
	assign w27709 = w27748 ^ w27706;
	assign w27753 = w27772 & w27803;
	assign w27747 = w27764 & w27812;
	assign w27746 = w27768 & w27809;
	assign w27712 = w27757 ^ w27746;
	assign w27708 = ~w27712;
	assign w27813 = w27708 ^ w27709;
	assign w44530 = w27747 ^ w27748;
	assign w27729 = w27753 ^ w44530;
	assign w27705 = w27729 ^ w27706;
	assign w49479 = w27704 ^ w27705;
	assign w27730 = w27754 ^ w27729;
	assign w49482 = w27730 ^ w27701;
	assign w27734 = w27762 ^ w27730;
	assign w27703 = w27761 ^ w27734;
	assign w49480 = w27702 ^ w27703;
	assign w27739 = w27763 ^ w27734;
	assign w27814 = w27739 ^ w27713;
	assign w49481 = w44531 ^ w27739;
	assign w27716 = w27720 ^ w44530;
	assign w27719 = w44532 ^ w27716;
	assign w27816 = w27718 ^ w27719;
	assign w27715 = w27711 ^ w27716;
	assign w27815 = w27714 ^ w27715;
	assign w45530 = ~w24600;
	assign w8495 = w45397 ^ w45530;
	assign w45535 = ~w24597;
	assign w45536 = ~w24598;
	assign w8468 = w45395 ^ w45536;
	assign w45537 = ~w24599;
	assign w8475 = w45396 ^ w45537;
	assign w45622 = ~w27814;
	assign w45623 = ~w27815;
	assign w45624 = ~w27816;
	assign w45629 = ~w27813;
	assign w45923 = ~w7974;
	assign w7762 = w45923 ^ w45261;
	assign w8044 = w7762 ^ w7763;
	assign w49122 = w8044 ^ w8036;
	assign w47243 = w49122 ^ w1701;
	assign w12847 = w47243 ^ w47241;
	assign w12937 = w47237 ^ w47243;
	assign w12849 = w47242 ^ w12847;
	assign w12922 = w47239 ^ w12849;
	assign w12918 = w12937 & w12922;
	assign w12924 = w12854 ^ w12849;
	assign w12916 = w12931 & w12924;
	assign w12852 = w12918 ^ w12848;
	assign w12925 = w47238 ^ w12849;
	assign w7898 = w45923 ^ w49260;
	assign w7919 = w45923 ^ w49243;
	assign w49136 = w7898 ^ w7899;
	assign w47229 = w49136 ^ w1715;
	assign w8191 = w47229 ^ w47235;
	assign w8189 = w47229 ^ w47234;
	assign w8172 = w8191 & w8176;
	assign w8190 = w47232 ^ w47229;
	assign w8169 = w8190 & w8179;
	assign w8105 = w8169 ^ w8103;
	assign w8182 = w8101 ^ w8190;
	assign w8102 = w47231 ^ w47229;
	assign w8185 = w8102 ^ w8108;
	assign w8064 = w8104 ^ w8102;
	assign w8180 = w8101 ^ w8064;
	assign w8167 = w8189 & w8180;
	assign w8170 = w8185 & w8178;
	assign w8177 = w8102 ^ w8192;
	assign w8168 = w8192 & w8177;
	assign w8077 = w8168 ^ w8169;
	assign w8124 = w8077 ^ w8078;
	assign w8183 = w8118 ^ w8185;
	assign w8106 = w8172 ^ w8102;
	assign w8186 = w8190 ^ w8118;
	assign w8175 = w8182 & w8186;
	assign w8107 = w8175 ^ w8104;
	assign w8111 = w8107 ^ w8105;
	assign w8116 = w47229 ^ w8111;
	assign w8181 = w47236 ^ w8182;
	assign w8174 = w8183 & w8181;
	assign w12930 = w47243 ^ w12934;
	assign w12917 = w12934 & w12930;
	assign w12864 = w47243 ^ w47242;
	assign w12929 = w12864 ^ w12931;
	assign w49125 = w7918 ^ w7919;
	assign w47240 = w49125 ^ w1704;
	assign w12936 = w47240 ^ w47237;
	assign w12932 = w12936 ^ w12864;
	assign w12915 = w12936 & w12925;
	assign w12851 = w12915 ^ w12849;
	assign w12928 = w12847 ^ w12936;
	assign w12921 = w12928 & w12932;
	assign w12927 = w47244 ^ w12928;
	assign w12920 = w12929 & w12927;
	assign w8125 = w8168 ^ w8174;
	assign w8166 = w8125 ^ w8116;
	assign w8123 = w8124 ^ w8106;
	assign w8165 = w8171 ^ w8123;
	assign w12850 = w47240 ^ w47238;
	assign w12810 = w12850 ^ w12848;
	assign w12926 = w12847 ^ w12810;
	assign w12913 = w12935 & w12926;
	assign w12809 = w12850 ^ w47239;
	assign w12933 = w47244 ^ w12809;
	assign w12919 = w47244 & w12933;
	assign w43798 = w8167 ^ w8173;
	assign w8079 = w8111 ^ w43798;
	assign w43799 = w8167 ^ w8170;
	assign w8120 = w8168 ^ w43799;
	assign w8076 = w8171 ^ w8120;
	assign w8158 = w47235 ^ w8076;
	assign w8080 = w8106 ^ w43799;
	assign w8164 = w8080 ^ w8105;
	assign w43908 = w12913 ^ w12919;
	assign w12863 = w43908 ^ w12848;
	assign w43909 = w12913 ^ w12916;
	assign w12826 = w12852 ^ w43909;
	assign w12910 = w12826 ^ w12851;
	assign w12938 = w47242 ^ w47240;
	assign w12923 = w12848 ^ w12938;
	assign w12914 = w12938 & w12923;
	assign w12866 = w12914 ^ w43909;
	assign w12823 = w12914 ^ w12915;
	assign w12822 = w12917 ^ w12866;
	assign w12870 = w12823 ^ w12824;
	assign w12904 = w47243 ^ w12822;
	assign w12869 = w12870 ^ w12852;
	assign w12911 = w12917 ^ w12869;
	assign w12871 = w12914 ^ w12920;
	assign w12909 = w12871 ^ w12863;
	assign w8122 = w47231 ^ w8079;
	assign w8162 = w8166 & w8165;
	assign w8161 = w8162 ^ w8164;
	assign w8157 = w8162 ^ w8122;
	assign w8156 = w8157 & w8158;
	assign w8075 = w8156 ^ w8120;
	assign w8074 = w8156 ^ w8173;
	assign w8069 = w8074 ^ w8170;
	assign w8154 = w8162 ^ w8156;
	assign w8153 = w8164 & w8154;
	assign w8151 = w8153 ^ w8161;
	assign w8155 = w8156 ^ w8164;
	assign w8132 = w8155 & w8187;
	assign w8141 = w8155 & w47236;
	assign w43802 = w8153 ^ w8171;
	assign w8145 = w43802 ^ w8123;
	assign w8143 = w8145 & w8182;
	assign w43801 = w8141 ^ w8143;
	assign w8112 = w47235 ^ w43802;
	assign w8152 = w8112 ^ w8075;
	assign w8142 = w8152 & w8181;
	assign w8134 = w8145 & w8186;
	assign w8133 = w8152 & w8183;
	assign w8117 = w43798 ^ w8102;
	assign w8163 = w8125 ^ w8117;
	assign w8160 = w8163 & w8161;
	assign w8068 = w8160 ^ w8116;
	assign w8071 = w8160 ^ w8172;
	assign w8067 = w8071 ^ w8107;
	assign w8070 = w47229 ^ w8067;
	assign w8066 = w47231 ^ w8067;
	assign w8147 = w8069 ^ w8070;
	assign w8128 = w8147 & w8190;
	assign w8137 = w8147 & w8179;
	assign w8159 = w8160 ^ w8122;
	assign w8129 = w8159 & w8185;
	assign w8138 = w8159 & w8178;
	assign w8150 = w8159 & w8151;
	assign w8073 = w8150 ^ w8174;
	assign w8115 = w8150 ^ w8125;
	assign w8149 = w8115 ^ w8117;
	assign w8139 = w8149 & w8188;
	assign w8082 = w8138 ^ w8139;
	assign w8130 = w8149 & w8184;
	assign w8100 = w8138 ^ w8130;
	assign w8146 = w8115 ^ w8068;
	assign w8131 = w8146 & w8191;
	assign w8140 = w8146 & w8176;
	assign w43800 = w8139 ^ w8140;
	assign w8098 = w8140 ^ w8131;
	assign w8065 = w8112 ^ w8073;
	assign w8072 = w8102 ^ w8065;
	assign w8148 = w8069 ^ w8072;
	assign w8126 = w8148 & w8189;
	assign w8144 = w8065 ^ w8066;
	assign w8127 = w8144 & w8192;
	assign w8092 = w8137 ^ w8126;
	assign w8136 = w8144 & w8177;
	assign w8135 = w8148 & w8180;
	assign w8113 = w8131 ^ w8135;
	assign w8121 = w8136 ^ w43800;
	assign w8097 = w8136 ^ w8139;
	assign w8088 = ~w8092;
	assign w8087 = w8132 ^ w8121;
	assign w8093 = w8136 ^ w8137;
	assign w8091 = ~w8113;
	assign w8081 = w8137 ^ w8121;
	assign w8090 = w8091 ^ w8129;
	assign w8086 = w8090 ^ w43801;
	assign w8089 = w8128 ^ w8086;
	assign w8193 = w8088 ^ w8089;
	assign w43523 = w8127 ^ w8128;
	assign w8109 = w8133 ^ w43523;
	assign w8085 = w8109 ^ w8086;
	assign w8096 = w8100 ^ w43523;
	assign w8099 = w43801 ^ w8096;
	assign w8196 = w8098 ^ w8099;
	assign w8084 = ~w8087;
	assign w8094 = ~w8097;
	assign w45201 = ~w8196;
	assign w8486 = w45201 ^ w45711;
	assign w8326 = w8488 ^ w8486;
	assign w8216 = w45201 ^ w45253;
	assign w8364 = w8486 ^ w8458;
	assign w49346 = w45253 ^ w8364;
	assign w47092 = w49346 ^ w1787;
	assign w8352 = w8486 ^ w8449;
	assign w49354 = w45401 ^ w8352;
	assign w47084 = w49354 ^ w1795;
	assign w45202 = ~w8193;
	assign w8464 = w45202 ^ w45716;
	assign w8360 = w8464 ^ w49477;
	assign w8342 = w8477 ^ w8464;
	assign w49359 = w45398 ^ w8342;
	assign w47079 = w49359 ^ w1800;
	assign w49351 = w8360 ^ w8361;
	assign w47087 = w49351 ^ w1792;
	assign w8330 = w8467 ^ w45202;
	assign w49368 = w8330 ^ w8331;
	assign w47070 = w49368 ^ w1809;
	assign w8095 = w8091 ^ w8096;
	assign w8195 = w8094 ^ w8095;
	assign w45204 = ~w8195;
	assign w8482 = w45204 ^ w45710;
	assign w8336 = w45204 ^ w12673;
	assign w49347 = w8537 ^ w8482;
	assign w49364 = w8335 ^ w8336;
	assign w47074 = w49364 ^ w1805;
	assign w8325 = w8484 ^ w8482;
	assign w8350 = w8489 ^ w8482;
	assign w47091 = w49347 ^ w1788;
	assign w8110 = w8134 ^ w8109;
	assign w49474 = w8110 ^ w8081;
	assign w8448 = w49474 ^ w49478;
	assign w8327 = w8448 ^ w45204;
	assign w49371 = w8326 ^ w8327;
	assign w8339 = w8448 ^ w45252;
	assign w8456 = w49470 ^ w49474;
	assign w8217 = w8456 ^ w49476;
	assign w8215 = w8456 ^ w45710;
	assign w8532 = w8215 ^ w8216;
	assign w49363 = w8532 ^ w8488;
	assign w47075 = w49363 ^ w1804;
	assign w8338 = w8489 ^ w8456;
	assign w8328 = w8489 ^ w8448;
	assign w49370 = w45201 ^ w8328;
	assign w8221 = ~w8456;
	assign w8219 = w8221 ^ w49477;
	assign w8114 = w8142 ^ w8110;
	assign w8119 = w8143 ^ w8114;
	assign w49473 = w43800 ^ w8119;
	assign w8194 = w8119 ^ w8093;
	assign w8469 = w49473 ^ w49477;
	assign w8318 = ~w49473;
	assign w8333 = w8318 ^ w49469;
	assign w49367 = w8332 ^ w8333;
	assign w47071 = w49367 ^ w1808;
	assign w8343 = w8345 ^ w8469;
	assign w8315 = w8473 ^ w8469;
	assign w49375 = w45202 ^ w8315;
	assign w47063 = w49375 ^ w1816;
	assign w47068 = w49370 ^ w1811;
	assign w49361 = w8339 ^ w8340;
	assign w47077 = w49361 ^ w1802;
	assign w33484 = w47079 ^ w47077;
	assign w17688 = w47075 ^ w47074;
	assign w8357 = w8467 ^ w8448;
	assign w49353 = w49470 ^ w8357;
	assign w47085 = w49353 ^ w1794;
	assign w17895 = w47085 ^ w47091;
	assign w17806 = w47087 ^ w47085;
	assign w47067 = w49371 ^ w1812;
	assign w8083 = w8141 ^ w8114;
	assign w49472 = w8082 ^ w8083;
	assign w8220 = w49472 ^ w8208;
	assign w8324 = w8448 ^ w49472;
	assign w8474 = w49472 ^ w49476;
	assign w8346 = w8337 ^ w8474;
	assign w8316 = w8319 ^ w8474;
	assign w8530 = w8219 ^ w8220;
	assign w49366 = w8530 ^ w8477;
	assign w47072 = w49366 ^ w1807;
	assign w17762 = w47074 ^ w47072;
	assign w17674 = w47072 ^ w47070;
	assign w17633 = w17674 ^ w47071;
	assign w49350 = w8535 ^ w8469;
	assign w47088 = w49350 ^ w1791;
	assign w17894 = w47088 ^ w47085;
	assign w8317 = w8448 ^ w8318;
	assign w49374 = w8316 ^ w8317;
	assign w47064 = w49374 ^ w1815;
	assign w49349 = w8536 ^ w8474;
	assign w47089 = w49349 ^ w1790;
	assign w17805 = w47091 ^ w47089;
	assign w45203 = ~w8194;
	assign w8466 = w45252 ^ w45203;
	assign w8329 = w8466 ^ w8449;
	assign w8314 = w8466 ^ w8464;
	assign w8358 = w8466 ^ w45717;
	assign w49352 = w8358 ^ w8359;
	assign w8313 = w49474 ^ w45203;
	assign w49377 = w8312 ^ w8313;
	assign w47061 = w49377 ^ w1818;
	assign w30536 = w47063 ^ w47061;
	assign w30624 = w47064 ^ w47061;
	assign w30625 = w47061 ^ w47067;
	assign w49369 = w49478 ^ w8329;
	assign w47069 = w49369 ^ w1810;
	assign w17759 = w47069 ^ w47074;
	assign w17672 = w47071 ^ w47069;
	assign w17761 = w47069 ^ w47075;
	assign w47086 = w49352 ^ w1793;
	assign w17812 = w47092 ^ w47086;
	assign w17892 = w47087 ^ w17812;
	assign w17888 = w47091 ^ w17892;
	assign w17875 = w17892 & w17888;
	assign w17889 = w17806 ^ w17812;
	assign w17634 = w17674 ^ w17672;
	assign w17747 = w17672 ^ w17762;
	assign w17738 = w17762 & w17747;
	assign w17760 = w47072 ^ w47069;
	assign w17756 = w17760 ^ w17688;
	assign w49376 = w45399 ^ w8314;
	assign w47062 = w49376 ^ w1817;
	assign w30538 = w47064 ^ w47062;
	assign w30542 = w47068 ^ w47062;
	assign w30619 = w30536 ^ w30542;
	assign w30622 = w47063 ^ w30542;
	assign w30618 = w47067 ^ w30622;
	assign w30498 = w30538 ^ w30536;
	assign w30497 = w30538 ^ w47063;
	assign w30621 = w47068 ^ w30497;
	assign w30607 = w47068 & w30621;
	assign w30605 = w30622 & w30618;
	assign w17808 = w47088 ^ w47086;
	assign w17768 = w17808 ^ w17806;
	assign w17884 = w17805 ^ w17768;
	assign w17767 = w17808 ^ w47087;
	assign w17891 = w47092 ^ w17767;
	assign w17877 = w47092 & w17891;
	assign w49362 = w45711 ^ w8338;
	assign w47076 = w49362 ^ w1803;
	assign w17757 = w47076 ^ w17633;
	assign w17678 = w47076 ^ w47070;
	assign w17758 = w47071 ^ w17678;
	assign w17754 = w47075 ^ w17758;
	assign w17755 = w17672 ^ w17678;
	assign w17743 = w47076 & w17757;
	assign w17741 = w17758 & w17754;
	assign w17753 = w17688 ^ w17755;
	assign w49360 = w45203 ^ w8341;
	assign w47078 = w49360 ^ w1801;
	assign w33490 = w47084 ^ w47078;
	assign w33567 = w33484 ^ w33490;
	assign w33570 = w47079 ^ w33490;
	assign w12853 = w12921 ^ w12850;
	assign w12857 = w12853 ^ w12851;
	assign w12825 = w12857 ^ w43908;
	assign w12868 = w47239 ^ w12825;
	assign w12862 = w47237 ^ w12857;
	assign w12912 = w12871 ^ w12862;
	assign w12908 = w12912 & w12911;
	assign w12903 = w12908 ^ w12868;
	assign w12902 = w12903 & w12904;
	assign w12900 = w12908 ^ w12902;
	assign w12821 = w12902 ^ w12866;
	assign w12820 = w12902 ^ w12919;
	assign w12899 = w12910 & w12900;
	assign w12815 = w12820 ^ w12916;
	assign w12901 = w12902 ^ w12910;
	assign w12887 = w12901 & w47244;
	assign w12878 = w12901 & w12933;
	assign w12907 = w12908 ^ w12910;
	assign w12897 = w12899 ^ w12907;
	assign w12906 = w12909 & w12907;
	assign w12905 = w12906 ^ w12868;
	assign w12884 = w12905 & w12924;
	assign w12875 = w12905 & w12931;
	assign w12817 = w12906 ^ w12918;
	assign w12813 = w12817 ^ w12853;
	assign w12812 = w47239 ^ w12813;
	assign w12896 = w12905 & w12897;
	assign w12819 = w12896 ^ w12920;
	assign w12861 = w12896 ^ w12871;
	assign w12895 = w12861 ^ w12863;
	assign w12885 = w12895 & w12934;
	assign w12828 = w12884 ^ w12885;
	assign w12876 = w12895 & w12930;
	assign w12846 = w12884 ^ w12876;
	assign w43913 = w12899 ^ w12917;
	assign w12891 = w43913 ^ w12869;
	assign w12889 = w12891 & w12928;
	assign w12880 = w12891 & w12932;
	assign w12858 = w47243 ^ w43913;
	assign w12811 = w12858 ^ w12819;
	assign w12890 = w12811 ^ w12812;
	assign w12873 = w12890 & w12938;
	assign w12882 = w12890 & w12923;
	assign w12843 = w12882 ^ w12885;
	assign w12840 = ~w12843;
	assign w12898 = w12858 ^ w12821;
	assign w12888 = w12898 & w12927;
	assign w12879 = w12898 & w12929;
	assign w12818 = w12848 ^ w12811;
	assign w12894 = w12815 ^ w12818;
	assign w12881 = w12894 & w12926;
	assign w12872 = w12894 & w12935;
	assign w43912 = w12887 ^ w12889;
	assign w12816 = w47237 ^ w12813;
	assign w12893 = w12815 ^ w12816;
	assign w12883 = w12893 & w12925;
	assign w12839 = w12882 ^ w12883;
	assign w12874 = w12893 & w12936;
	assign w12838 = w12883 ^ w12872;
	assign w12834 = ~w12838;
	assign w43910 = w12873 ^ w12874;
	assign w12855 = w12879 ^ w43910;
	assign w12856 = w12880 ^ w12855;
	assign w12860 = w12888 ^ w12856;
	assign w12865 = w12889 ^ w12860;
	assign w12940 = w12865 ^ w12839;
	assign w8273 = w45626 ^ w12940;
	assign w8301 = w12940 ^ w45629;
	assign w49488 = ~w12940;
	assign w8476 = w45622 ^ w49488;
	assign w12829 = w12887 ^ w12860;
	assign w49485 = w12828 ^ w12829;
	assign w8498 = w49480 ^ w49485;
	assign w8265 = ~w8498;
	assign w12842 = w12846 ^ w43910;
	assign w12845 = w43912 ^ w12842;
	assign w12814 = w12906 ^ w12862;
	assign w12892 = w12861 ^ w12814;
	assign w12886 = w12892 & w12922;
	assign w12877 = w12892 & w12937;
	assign w12859 = w12877 ^ w12881;
	assign w12844 = w12886 ^ w12877;
	assign w43911 = w12885 ^ w12886;
	assign w12867 = w12882 ^ w43911;
	assign w12833 = w12878 ^ w12867;
	assign w12830 = ~w12833;
	assign w12827 = w12883 ^ w12867;
	assign w49489 = w12856 ^ w12827;
	assign w8298 = w49489 ^ w45622;
	assign w8454 = w49489 ^ w49493;
	assign w8235 = ~w8454;
	assign w8450 = w49482 ^ w49489;
	assign w49486 = w43911 ^ w12865;
	assign w8278 = w49492 ^ w49486;
	assign w8229 = w49486 ^ w49480;
	assign w8490 = w49481 ^ w49486;
	assign w8262 = ~w8490;
	assign w12942 = w12844 ^ w12845;
	assign w12837 = ~w12859;
	assign w12841 = w12837 ^ w12842;
	assign w12941 = w12840 ^ w12841;
	assign w8280 = w45627 ^ w12941;
	assign w12836 = w12837 ^ w12875;
	assign w12832 = w12836 ^ w43912;
	assign w12835 = w12874 ^ w12832;
	assign w12939 = w12834 ^ w12835;
	assign w8306 = w12939 ^ w49481;
	assign w12831 = w12855 ^ w12832;
	assign w49484 = w12830 ^ w12831;
	assign w8234 = ~w49484;
	assign w8505 = w49479 ^ w49484;
	assign w49483 = ~w12941;
	assign w8512 = w45623 ^ w49483;
	assign w8233 = w49490 ^ w8234;
	assign w49487 = ~w12939;
	assign w8483 = w45629 ^ w49487;
	assign w8281 = ~w8505;
	assign w8275 = w45633 ^ w12939;
	assign w8227 = ~w49485;
	assign w8226 = w8227 ^ w49479;
	assign w8237 = w49491 ^ w8227;
	assign w45254 = ~w12942;
	assign w8231 = w45628 ^ w45254;
	assign w8513 = w45624 ^ w45254;
	assign w8282 = w8513 ^ w8454;
	assign w8309 = w8234 ^ w45623;
	assign w49471 = w8084 ^ w8085;
	assign w8218 = w49471 ^ w49467;
	assign w8531 = w8217 ^ w8218;
	assign w8479 = w49471 ^ w49475;
	assign w8348 = w8488 ^ w8479;
	assign w49372 = w49471 ^ w8325;
	assign w47066 = w49372 ^ w1813;
	assign w30552 = w47067 ^ w47066;
	assign w30617 = w30552 ^ w30619;
	assign w30620 = w30624 ^ w30552;
	assign w30626 = w47066 ^ w47064;
	assign w30611 = w30536 ^ w30626;
	assign w30623 = w47061 ^ w47066;
	assign w30602 = w30626 & w30611;
	assign w8362 = w8479 ^ w45710;
	assign w49348 = w8362 ^ w8363;
	assign w47090 = w49348 ^ w1789;
	assign w17893 = w47085 ^ w47090;
	assign w17871 = w17893 & w17884;
	assign w17782 = w47089 ^ w47090;
	assign w17807 = w47090 ^ w17805;
	assign w17822 = w47091 ^ w47090;
	assign w17890 = w17894 ^ w17822;
	assign w17882 = w17812 ^ w17807;
	assign w17874 = w17889 & w17882;
	assign w17880 = w47087 ^ w17807;
	assign w17876 = w17895 & w17880;
	assign w17810 = w17876 ^ w17806;
	assign w17883 = w47086 ^ w17807;
	assign w17873 = w17894 & w17883;
	assign w17896 = w47090 ^ w47088;
	assign w17881 = w17806 ^ w17896;
	assign w17872 = w17896 & w17881;
	assign w17781 = w17872 ^ w17873;
	assign w17828 = w17781 ^ w17782;
	assign w17827 = w17828 ^ w17810;
	assign w17869 = w17875 ^ w17827;
	assign w49356 = w49462 ^ w8348;
	assign w47082 = w49356 ^ w1797;
	assign w33571 = w47077 ^ w47082;
	assign w44116 = w17871 ^ w17874;
	assign w17824 = w17872 ^ w44116;
	assign w17780 = w17875 ^ w17824;
	assign w17862 = w47091 ^ w17780;
	assign w17784 = w17810 ^ w44116;
	assign w49365 = w8531 ^ w8481;
	assign w47073 = w49365 ^ w1806;
	assign w17671 = w47075 ^ w47073;
	assign w17750 = w17671 ^ w17634;
	assign w17737 = w17759 & w17750;
	assign w17752 = w17671 ^ w17760;
	assign w17751 = w47076 ^ w17752;
	assign w17744 = w17753 & w17751;
	assign w17648 = w47073 ^ w47074;
	assign w17673 = w47074 ^ w17671;
	assign w17749 = w47070 ^ w17673;
	assign w17739 = w17760 & w17749;
	assign w17647 = w17738 ^ w17739;
	assign w17694 = w17647 ^ w17648;
	assign w17746 = w47071 ^ w17673;
	assign w17742 = w17761 & w17746;
	assign w17676 = w17742 ^ w17672;
	assign w17675 = w17739 ^ w17673;
	assign w17693 = w17694 ^ w17676;
	assign w17735 = w17741 ^ w17693;
	assign w17748 = w17678 ^ w17673;
	assign w17740 = w17755 & w17748;
	assign w17745 = w17752 & w17756;
	assign w17677 = w17745 ^ w17674;
	assign w17681 = w17677 ^ w17675;
	assign w17686 = w47069 ^ w17681;
	assign w44109 = w17737 ^ w17740;
	assign w17650 = w17676 ^ w44109;
	assign w17734 = w17650 ^ w17675;
	assign w44112 = w17737 ^ w17743;
	assign w17649 = w17681 ^ w44112;
	assign w17692 = w47071 ^ w17649;
	assign w17687 = w44112 ^ w17672;
	assign w17690 = w17738 ^ w44109;
	assign w17646 = w17741 ^ w17690;
	assign w17728 = w47075 ^ w17646;
	assign w8323 = w8481 ^ w8479;
	assign w49373 = w8323 ^ w8324;
	assign w47065 = w49373 ^ w1814;
	assign w30535 = w47067 ^ w47065;
	assign w30537 = w47066 ^ w30535;
	assign w30613 = w47062 ^ w30537;
	assign w30610 = w47063 ^ w30537;
	assign w30612 = w30542 ^ w30537;
	assign w30616 = w30535 ^ w30624;
	assign w30615 = w47068 ^ w30616;
	assign w30512 = w47065 ^ w47066;
	assign w30614 = w30535 ^ w30498;
	assign w30609 = w30616 & w30620;
	assign w30541 = w30609 ^ w30538;
	assign w30608 = w30617 & w30615;
	assign w30559 = w30602 ^ w30608;
	assign w30606 = w30625 & w30610;
	assign w30540 = w30606 ^ w30536;
	assign w30604 = w30619 & w30612;
	assign w30603 = w30624 & w30613;
	assign w30539 = w30603 ^ w30537;
	assign w30545 = w30541 ^ w30539;
	assign w30550 = w47061 ^ w30545;
	assign w30600 = w30559 ^ w30550;
	assign w30511 = w30602 ^ w30603;
	assign w30558 = w30511 ^ w30512;
	assign w30557 = w30558 ^ w30540;
	assign w30599 = w30605 ^ w30557;
	assign w30601 = w30623 & w30614;
	assign w30596 = w30600 & w30599;
	assign w17887 = w17822 ^ w17889;
	assign w44649 = w30601 ^ w30607;
	assign w30551 = w44649 ^ w30536;
	assign w30597 = w30559 ^ w30551;
	assign w30513 = w30545 ^ w44649;
	assign w30556 = w47063 ^ w30513;
	assign w30591 = w30596 ^ w30556;
	assign w44650 = w30601 ^ w30604;
	assign w30554 = w30602 ^ w44650;
	assign w30510 = w30605 ^ w30554;
	assign w30592 = w47067 ^ w30510;
	assign w30590 = w30591 & w30592;
	assign w30509 = w30590 ^ w30554;
	assign w30508 = w30590 ^ w30607;
	assign w30503 = w30508 ^ w30604;
	assign w30588 = w30596 ^ w30590;
	assign w30514 = w30540 ^ w44650;
	assign w30598 = w30514 ^ w30539;
	assign w30589 = w30590 ^ w30598;
	assign w30595 = w30596 ^ w30598;
	assign w30594 = w30597 & w30595;
	assign w30593 = w30594 ^ w30556;
	assign w30505 = w30594 ^ w30606;
	assign w30501 = w30505 ^ w30541;
	assign w30504 = w47061 ^ w30501;
	assign w30581 = w30503 ^ w30504;
	assign w30502 = w30594 ^ w30550;
	assign w30500 = w47063 ^ w30501;
	assign w30587 = w30598 & w30588;
	assign w30585 = w30587 ^ w30595;
	assign w30584 = w30593 & w30585;
	assign w30549 = w30584 ^ w30559;
	assign w30583 = w30549 ^ w30551;
	assign w30507 = w30584 ^ w30608;
	assign w30580 = w30549 ^ w30502;
	assign w30575 = w30589 & w47068;
	assign w30574 = w30580 & w30610;
	assign w30573 = w30583 & w30622;
	assign w30572 = w30593 & w30612;
	assign w30516 = w30572 ^ w30573;
	assign w30571 = w30581 & w30613;
	assign w30566 = w30589 & w30621;
	assign w30565 = w30580 & w30625;
	assign w30532 = w30574 ^ w30565;
	assign w30564 = w30583 & w30618;
	assign w30534 = w30572 ^ w30564;
	assign w30563 = w30593 & w30619;
	assign w30562 = w30581 & w30624;
	assign w44651 = w30573 ^ w30574;
	assign w44653 = w30587 ^ w30605;
	assign w30546 = w47067 ^ w44653;
	assign w30586 = w30546 ^ w30509;
	assign w30567 = w30586 & w30617;
	assign w30576 = w30586 & w30615;
	assign w30499 = w30546 ^ w30507;
	assign w30506 = w30536 ^ w30499;
	assign w30582 = w30503 ^ w30506;
	assign w30569 = w30582 & w30614;
	assign w30547 = w30565 ^ w30569;
	assign w30525 = ~w30547;
	assign w30524 = w30525 ^ w30563;
	assign w30578 = w30499 ^ w30500;
	assign w30561 = w30578 & w30626;
	assign w30560 = w30582 & w30623;
	assign w30526 = w30571 ^ w30560;
	assign w30522 = ~w30526;
	assign w43584 = w30561 ^ w30562;
	assign w30530 = w30534 ^ w43584;
	assign w30529 = w30525 ^ w30530;
	assign w30543 = w30567 ^ w43584;
	assign w30570 = w30578 & w30611;
	assign w30527 = w30570 ^ w30571;
	assign w30555 = w30570 ^ w44651;
	assign w30521 = w30566 ^ w30555;
	assign w30518 = ~w30521;
	assign w30515 = w30571 ^ w30555;
	assign w30531 = w30570 ^ w30573;
	assign w30528 = ~w30531;
	assign w30629 = w30528 ^ w30529;
	assign w30579 = w44653 ^ w30557;
	assign w30577 = w30579 & w30616;
	assign w30568 = w30579 & w30620;
	assign w30544 = w30568 ^ w30543;
	assign w30548 = w30576 ^ w30544;
	assign w30553 = w30577 ^ w30548;
	assign w49678 = w44651 ^ w30553;
	assign w30628 = w30553 ^ w30527;
	assign w30517 = w30575 ^ w30548;
	assign w49677 = w30516 ^ w30517;
	assign w49679 = w30544 ^ w30515;
	assign w44652 = w30575 ^ w30577;
	assign w30533 = w44652 ^ w30530;
	assign w30630 = w30532 ^ w30533;
	assign w30520 = w30524 ^ w44652;
	assign w30523 = w30562 ^ w30520;
	assign w30627 = w30522 ^ w30523;
	assign w30519 = w30543 ^ w30520;
	assign w49676 = w30518 ^ w30519;
	assign w17809 = w17873 ^ w17807;
	assign w17868 = w17784 ^ w17809;
	assign w45698 = ~w30630;
	assign w45703 = ~w30627;
	assign w45704 = ~w30628;
	assign w45705 = ~w30629;
	assign w44115 = w17871 ^ w17877;
	assign w17821 = w44115 ^ w17806;
	assign w45891 = ~w8450;
	assign w8295 = w45891 ^ w45623;
	assign w8289 = w45891 ^ w49481;
	assign w8291 = w45891 ^ w49480;
	assign w17695 = w17738 ^ w17744;
	assign w17733 = w17695 ^ w17687;
	assign w17736 = w17695 ^ w17686;
	assign w17732 = w17736 & w17735;
	assign w17731 = w17732 ^ w17734;
	assign w17730 = w17733 & w17731;
	assign w17638 = w17730 ^ w17686;
	assign w17641 = w17730 ^ w17742;
	assign w17637 = w17641 ^ w17677;
	assign w17640 = w47069 ^ w17637;
	assign w17729 = w17730 ^ w17692;
	assign w17708 = w17729 & w17748;
	assign w17699 = w17729 & w17755;
	assign w17636 = w47071 ^ w17637;
	assign w17727 = w17732 ^ w17692;
	assign w17726 = w17727 & w17728;
	assign w17644 = w17726 ^ w17743;
	assign w17639 = w17644 ^ w17740;
	assign w17645 = w17726 ^ w17690;
	assign w17717 = w17639 ^ w17640;
	assign w17707 = w17717 & w17749;
	assign w17698 = w17717 & w17760;
	assign w17725 = w17726 ^ w17734;
	assign w17724 = w17732 ^ w17726;
	assign w17723 = w17734 & w17724;
	assign w17721 = w17723 ^ w17731;
	assign w17720 = w17729 & w17721;
	assign w17643 = w17720 ^ w17744;
	assign w17711 = w17725 & w47076;
	assign w17702 = w17725 & w17757;
	assign w44111 = w17723 ^ w17741;
	assign w17715 = w44111 ^ w17693;
	assign w17713 = w17715 & w17752;
	assign w44114 = w17711 ^ w17713;
	assign w17704 = w17715 & w17756;
	assign w17682 = w47075 ^ w44111;
	assign w17722 = w17682 ^ w17645;
	assign w17635 = w17682 ^ w17643;
	assign w17642 = w17672 ^ w17635;
	assign w17718 = w17639 ^ w17642;
	assign w17696 = w17718 & w17759;
	assign w17662 = w17707 ^ w17696;
	assign w17658 = ~w17662;
	assign w17705 = w17718 & w17750;
	assign w17714 = w17635 ^ w17636;
	assign w17706 = w17714 & w17747;
	assign w17663 = w17706 ^ w17707;
	assign w17697 = w17714 & w17762;
	assign w17712 = w17722 & w17751;
	assign w17703 = w17722 & w17753;
	assign w44110 = w17697 ^ w17698;
	assign w17679 = w17703 ^ w44110;
	assign w17680 = w17704 ^ w17679;
	assign w17684 = w17712 ^ w17680;
	assign w17653 = w17711 ^ w17684;
	assign w17689 = w17713 ^ w17684;
	assign w17764 = w17689 ^ w17663;
	assign w45385 = ~w17764;
	assign w17685 = w17720 ^ w17695;
	assign w17716 = w17685 ^ w17638;
	assign w17719 = w17685 ^ w17687;
	assign w17709 = w17719 & w17758;
	assign w17667 = w17706 ^ w17709;
	assign w17664 = ~w17667;
	assign w17700 = w17719 & w17754;
	assign w17670 = w17708 ^ w17700;
	assign w17652 = w17708 ^ w17709;
	assign w17710 = w17716 & w17746;
	assign w17701 = w17716 & w17761;
	assign w17668 = w17710 ^ w17701;
	assign w17683 = w17701 ^ w17705;
	assign w49692 = w17652 ^ w17653;
	assign w17666 = w17670 ^ w44110;
	assign w17669 = w44114 ^ w17666;
	assign w17766 = w17668 ^ w17669;
	assign w17661 = ~w17683;
	assign w17660 = w17661 ^ w17699;
	assign w17656 = w17660 ^ w44114;
	assign w17659 = w17698 ^ w17656;
	assign w17763 = w17658 ^ w17659;
	assign w17655 = w17679 ^ w17656;
	assign w44113 = w17709 ^ w17710;
	assign w49693 = w44113 ^ w17689;
	assign w17691 = w17706 ^ w44113;
	assign w17657 = w17702 ^ w17691;
	assign w17654 = ~w17657;
	assign w17651 = w17707 ^ w17691;
	assign w49694 = w17680 ^ w17651;
	assign w49691 = w17654 ^ w17655;
	assign w45379 = ~w17766;
	assign w45384 = ~w17763;
	assign w17665 = w17661 ^ w17666;
	assign w17765 = w17664 ^ w17665;
	assign w45378 = ~w17765;
	assign w17886 = w17805 ^ w17894;
	assign w17879 = w17886 & w17890;
	assign w17811 = w17879 ^ w17808;
	assign w17815 = w17811 ^ w17809;
	assign w17783 = w17815 ^ w44115;
	assign w17826 = w47087 ^ w17783;
	assign w17820 = w47085 ^ w17815;
	assign w17885 = w47092 ^ w17886;
	assign w17878 = w17887 & w17885;
	assign w17829 = w17872 ^ w17878;
	assign w17870 = w17829 ^ w17820;
	assign w17866 = w17870 & w17869;
	assign w17861 = w17866 ^ w17826;
	assign w17860 = w17861 & w17862;
	assign w17778 = w17860 ^ w17877;
	assign w17773 = w17778 ^ w17874;
	assign w17859 = w17860 ^ w17868;
	assign w17845 = w17859 & w47092;
	assign w17836 = w17859 & w17891;
	assign w17858 = w17866 ^ w17860;
	assign w17857 = w17868 & w17858;
	assign w17865 = w17866 ^ w17868;
	assign w17855 = w17857 ^ w17865;
	assign w17867 = w17829 ^ w17821;
	assign w17864 = w17867 & w17865;
	assign w17775 = w17864 ^ w17876;
	assign w17771 = w17775 ^ w17811;
	assign w17770 = w47087 ^ w17771;
	assign w17774 = w47085 ^ w17771;
	assign w17863 = w17864 ^ w17826;
	assign w17854 = w17863 & w17855;
	assign w17833 = w17863 & w17889;
	assign w17842 = w17863 & w17882;
	assign w17777 = w17854 ^ w17878;
	assign w17819 = w17854 ^ w17829;
	assign w17853 = w17819 ^ w17821;
	assign w17843 = w17853 & w17892;
	assign w17834 = w17853 & w17888;
	assign w17804 = w17842 ^ w17834;
	assign w17786 = w17842 ^ w17843;
	assign w17851 = w17773 ^ w17774;
	assign w17832 = w17851 & w17894;
	assign w17841 = w17851 & w17883;
	assign w17772 = w17864 ^ w17820;
	assign w17850 = w17819 ^ w17772;
	assign w17844 = w17850 & w17880;
	assign w17835 = w17850 & w17895;
	assign w17802 = w17844 ^ w17835;
	assign w44117 = w17843 ^ w17844;
	assign w44119 = w17857 ^ w17875;
	assign w17816 = w47091 ^ w44119;
	assign w17769 = w17816 ^ w17777;
	assign w17848 = w17769 ^ w17770;
	assign w17840 = w17848 & w17881;
	assign w17797 = w17840 ^ w17841;
	assign w17831 = w17848 & w17896;
	assign w17825 = w17840 ^ w44117;
	assign w17791 = w17836 ^ w17825;
	assign w17785 = w17841 ^ w17825;
	assign w17788 = ~w17791;
	assign w43548 = w17831 ^ w17832;
	assign w17800 = w17804 ^ w43548;
	assign w17776 = w17806 ^ w17769;
	assign w17852 = w17773 ^ w17776;
	assign w17839 = w17852 & w17884;
	assign w17830 = w17852 & w17893;
	assign w17796 = w17841 ^ w17830;
	assign w17792 = ~w17796;
	assign w17817 = w17835 ^ w17839;
	assign w17795 = ~w17817;
	assign w17799 = w17795 ^ w17800;
	assign w17794 = w17795 ^ w17833;
	assign w17801 = w17840 ^ w17843;
	assign w17798 = ~w17801;
	assign w17899 = w17798 ^ w17799;
	assign w17849 = w44119 ^ w17827;
	assign w17847 = w17849 & w17886;
	assign w17838 = w17849 & w17890;
	assign w44118 = w17845 ^ w17847;
	assign w17803 = w44118 ^ w17800;
	assign w17900 = w17802 ^ w17803;
	assign w17790 = w17794 ^ w44118;
	assign w17793 = w17832 ^ w17790;
	assign w17897 = w17792 ^ w17793;
	assign w45382 = ~w17899;
	assign w45383 = ~w17900;
	assign w45388 = ~w17897;
	assign w17779 = w17860 ^ w17824;
	assign w17856 = w17816 ^ w17779;
	assign w17846 = w17856 & w17885;
	assign w17837 = w17856 & w17887;
	assign w17813 = w17837 ^ w43548;
	assign w17789 = w17813 ^ w17790;
	assign w17814 = w17838 ^ w17813;
	assign w49646 = w17814 ^ w17785;
	assign w49643 = w17788 ^ w17789;
	assign w17818 = w17846 ^ w17814;
	assign w17787 = w17845 ^ w17818;
	assign w49644 = w17786 ^ w17787;
	assign w17823 = w17847 ^ w17818;
	assign w17898 = w17823 ^ w17797;
	assign w49645 = w44117 ^ w17823;
	assign w45389 = ~w17898;
	assign w8223 = w12941 ^ w45624;
	assign w45924 = ~w7973;
	assign w7768 = w45924 ^ w49256;
	assign w8041 = w7768 ^ w7769;
	assign w7805 = w45924 ^ w45634;
	assign w49140 = w8041 ^ w8038;
	assign w47225 = w49140 ^ w1719;
	assign w24639 = w47227 ^ w47225;
	assign w24641 = w47226 ^ w24639;
	assign w24717 = w47222 ^ w24641;
	assign w24714 = w47223 ^ w24641;
	assign w24716 = w24646 ^ w24641;
	assign w24616 = w47225 ^ w47226;
	assign w24710 = w24729 & w24714;
	assign w24644 = w24710 ^ w24640;
	assign w24708 = w24723 & w24716;
	assign w7892 = w45924 ^ w49254;
	assign w49141 = w7891 ^ w7892;
	assign w47224 = w49141 ^ w1720;
	assign w24642 = w47224 ^ w47222;
	assign w24728 = w47224 ^ w47221;
	assign w24724 = w24728 ^ w24656;
	assign w24720 = w24639 ^ w24728;
	assign w24719 = w47228 ^ w24720;
	assign w24730 = w47226 ^ w47224;
	assign w24715 = w24640 ^ w24730;
	assign w24602 = w24642 ^ w24640;
	assign w24718 = w24639 ^ w24602;
	assign w24601 = w24642 ^ w47223;
	assign w24725 = w47228 ^ w24601;
	assign w24713 = w24720 & w24724;
	assign w24645 = w24713 ^ w24642;
	assign w24712 = w24721 & w24719;
	assign w24711 = w47228 & w24725;
	assign w24707 = w24728 & w24717;
	assign w24643 = w24707 ^ w24641;
	assign w24649 = w24645 ^ w24643;
	assign w24654 = w47221 ^ w24649;
	assign w24706 = w24730 & w24715;
	assign w24663 = w24706 ^ w24712;
	assign w24704 = w24663 ^ w24654;
	assign w24615 = w24706 ^ w24707;
	assign w24662 = w24615 ^ w24616;
	assign w24661 = w24662 ^ w24644;
	assign w24703 = w24709 ^ w24661;
	assign w24705 = w24727 & w24718;
	assign w24700 = w24704 & w24703;
	assign w49120 = w7805 ^ w7806;
	assign w44402 = w24705 ^ w24708;
	assign w24618 = w24644 ^ w44402;
	assign w24702 = w24618 ^ w24643;
	assign w24699 = w24700 ^ w24702;
	assign w24658 = w24706 ^ w44402;
	assign w24614 = w24709 ^ w24658;
	assign w24696 = w47227 ^ w24614;
	assign w44405 = w24705 ^ w24711;
	assign w24617 = w24649 ^ w44405;
	assign w24660 = w47223 ^ w24617;
	assign w24695 = w24700 ^ w24660;
	assign w24694 = w24695 & w24696;
	assign w24692 = w24700 ^ w24694;
	assign w24613 = w24694 ^ w24658;
	assign w24612 = w24694 ^ w24711;
	assign w24607 = w24612 ^ w24708;
	assign w24691 = w24702 & w24692;
	assign w24689 = w24691 ^ w24699;
	assign w44404 = w24691 ^ w24709;
	assign w24683 = w44404 ^ w24661;
	assign w24672 = w24683 & w24724;
	assign w24681 = w24683 & w24720;
	assign w24650 = w47227 ^ w44404;
	assign w24690 = w24650 ^ w24613;
	assign w24680 = w24690 & w24719;
	assign w24671 = w24690 & w24721;
	assign w24693 = w24694 ^ w24702;
	assign w24679 = w24693 & w47228;
	assign w24670 = w24693 & w24725;
	assign w24655 = w44405 ^ w24640;
	assign w24701 = w24663 ^ w24655;
	assign w24698 = w24701 & w24699;
	assign w24697 = w24698 ^ w24660;
	assign w24609 = w24698 ^ w24710;
	assign w24605 = w24609 ^ w24645;
	assign w24608 = w47221 ^ w24605;
	assign w24685 = w24607 ^ w24608;
	assign w24606 = w24698 ^ w24654;
	assign w24604 = w47223 ^ w24605;
	assign w24688 = w24697 & w24689;
	assign w24653 = w24688 ^ w24663;
	assign w24687 = w24653 ^ w24655;
	assign w24611 = w24688 ^ w24712;
	assign w24603 = w24650 ^ w24611;
	assign w24610 = w24640 ^ w24603;
	assign w24686 = w24607 ^ w24610;
	assign w24684 = w24653 ^ w24606;
	assign w24682 = w24603 ^ w24604;
	assign w24678 = w24684 & w24714;
	assign w24677 = w24687 & w24726;
	assign w24676 = w24697 & w24716;
	assign w24620 = w24676 ^ w24677;
	assign w24675 = w24685 & w24717;
	assign w24674 = w24682 & w24715;
	assign w24635 = w24674 ^ w24677;
	assign w24632 = ~w24635;
	assign w24631 = w24674 ^ w24675;
	assign w24673 = w24686 & w24718;
	assign w24669 = w24684 & w24729;
	assign w24651 = w24669 ^ w24673;
	assign w24636 = w24678 ^ w24669;
	assign w24629 = ~w24651;
	assign w24668 = w24687 & w24722;
	assign w24638 = w24676 ^ w24668;
	assign w24667 = w24697 & w24723;
	assign w24628 = w24629 ^ w24667;
	assign w24666 = w24685 & w24728;
	assign w24665 = w24682 & w24730;
	assign w24664 = w24686 & w24727;
	assign w24630 = w24675 ^ w24664;
	assign w24626 = ~w24630;
	assign w44403 = w24665 ^ w24666;
	assign w24647 = w24671 ^ w44403;
	assign w24648 = w24672 ^ w24647;
	assign w24652 = w24680 ^ w24648;
	assign w24621 = w24679 ^ w24652;
	assign w49458 = w24620 ^ w24621;
	assign w8506 = w49454 ^ w49458;
	assign w49325 = w8521 ^ w8506;
	assign w47113 = w49325 ^ w1830;
	assign w8371 = w8507 ^ w8506;
	assign w8369 = ~w8371;
	assign w8386 = w8387 ^ w49458;
	assign w49333 = w8385 ^ w8386;
	assign w47105 = w49333 ^ w1838;
	assign w8202 = w49458 ^ w49448;
	assign w24657 = w24681 ^ w24652;
	assign w24732 = w24657 ^ w24631;
	assign w49460 = ~w24732;
	assign w8496 = w45391 ^ w49460;
	assign w8394 = w8504 ^ w8496;
	assign w8303 = w8496 ^ w45402;
	assign w49328 = w45403 ^ w8394;
	assign w47110 = w49328 ^ w1833;
	assign w8378 = w8502 ^ w24732;
	assign w49336 = w8378 ^ w8379;
	assign w47102 = w49336 ^ w1841;
	assign w8284 = w24732 ^ w49451;
	assign w24634 = w24638 ^ w44403;
	assign w24633 = w24629 ^ w24634;
	assign w24733 = w24632 ^ w24633;
	assign w44406 = w24677 ^ w24678;
	assign w49459 = w44406 ^ w24657;
	assign w8503 = w49455 ^ w49459;
	assign w8238 = w8453 ^ w49459;
	assign w8396 = w8398 ^ w8503;
	assign w8368 = w8504 ^ w8503;
	assign w49343 = w45390 ^ w8368;
	assign w47095 = w49343 ^ w1848;
	assign w24659 = w24674 ^ w44406;
	assign w24625 = w24670 ^ w24659;
	assign w24622 = ~w24625;
	assign w24619 = w24675 ^ w24659;
	assign w49461 = w24648 ^ w24619;
	assign w8451 = w49456 ^ w49461;
	assign w8459 = w49445 ^ w49461;
	assign w8444 = w8492 ^ w8459;
	assign w8375 = w8492 ^ w8451;
	assign w49338 = w45405 ^ w8375;
	assign w47100 = w49338 ^ w1843;
	assign w8201 = w8459 ^ w49443;
	assign w8538 = w8201 ^ w8202;
	assign w49318 = w8538 ^ w8503;
	assign w8393 = w8502 ^ w8451;
	assign w49329 = w49445 ^ w8393;
	assign w47109 = w49329 ^ w1834;
	assign w47120 = w49318 ^ w1823;
	assign w8355 = ~w8459;
	assign w8354 = w8355 ^ w49447;
	assign w44407 = w24679 ^ w24681;
	assign w24637 = w44407 ^ w24634;
	assign w24734 = w24636 ^ w24637;
	assign w24624 = w24628 ^ w44407;
	assign w24627 = w24666 ^ w24624;
	assign w24731 = w24626 ^ w24627;
	assign w24623 = w24647 ^ w24624;
	assign w49457 = w24622 ^ w24623;
	assign w8494 = w49442 ^ w49457;
	assign w8388 = w8494 ^ w8493;
	assign w49332 = w49446 ^ w8388;
	assign w47106 = w49332 ^ w1837;
	assign w27564 = w47105 ^ w47106;
	assign w8356 = ~w8494;
	assign w8425 = w8356 ^ w45779;
	assign w49324 = w8425 ^ w8426;
	assign w47114 = w49324 ^ w1829;
	assign w12422 = w47113 ^ w47114;
	assign w12533 = w47109 ^ w47114;
	assign w8353 = w8506 ^ w8356;
	assign w49317 = w8353 ^ w8354;
	assign w47121 = w49317 ^ w1822;
	assign w8365 = w8496 ^ w8452;
	assign w49345 = w49456 ^ w8365;
	assign w47093 = w49345 ^ w1850;
	assign w30670 = w47095 ^ w47093;
	assign w8523 = w8238 ^ w8239;
	assign w49334 = w8523 ^ w8507;
	assign w47104 = w49334 ^ w1839;
	assign w27590 = w47104 ^ w47102;
	assign w27678 = w47106 ^ w47104;
	assign w47245 = w49120 ^ w1699;
	assign w24774 = w47247 ^ w47245;
	assign w24849 = w24774 ^ w24864;
	assign w24862 = w47248 ^ w47245;
	assign w24858 = w24862 ^ w24790;
	assign w24857 = w24774 ^ w24780;
	assign w24855 = w24790 ^ w24857;
	assign w24854 = w24773 ^ w24862;
	assign w24853 = w47252 ^ w24854;
	assign w24736 = w24776 ^ w24774;
	assign w24852 = w24773 ^ w24736;
	assign w24863 = w47245 ^ w47251;
	assign w24861 = w47245 ^ w47250;
	assign w24847 = w24854 & w24858;
	assign w24779 = w24847 ^ w24776;
	assign w24846 = w24855 & w24853;
	assign w24844 = w24863 & w24848;
	assign w24778 = w24844 ^ w24774;
	assign w24842 = w24857 & w24850;
	assign w24841 = w24862 & w24851;
	assign w24777 = w24841 ^ w24775;
	assign w24783 = w24779 ^ w24777;
	assign w24788 = w47245 ^ w24783;
	assign w24840 = w24864 & w24849;
	assign w24797 = w24840 ^ w24846;
	assign w24838 = w24797 ^ w24788;
	assign w24749 = w24840 ^ w24841;
	assign w24796 = w24749 ^ w24750;
	assign w24795 = w24796 ^ w24778;
	assign w24837 = w24843 ^ w24795;
	assign w24839 = w24861 & w24852;
	assign w24834 = w24838 & w24837;
	assign w44408 = w24839 ^ w24845;
	assign w24751 = w24783 ^ w44408;
	assign w24794 = w47247 ^ w24751;
	assign w24829 = w24834 ^ w24794;
	assign w24789 = w44408 ^ w24774;
	assign w24835 = w24797 ^ w24789;
	assign w44409 = w24839 ^ w24842;
	assign w24792 = w24840 ^ w44409;
	assign w24748 = w24843 ^ w24792;
	assign w24830 = w47251 ^ w24748;
	assign w24828 = w24829 & w24830;
	assign w24747 = w24828 ^ w24792;
	assign w24826 = w24834 ^ w24828;
	assign w24746 = w24828 ^ w24845;
	assign w24741 = w24746 ^ w24842;
	assign w24752 = w24778 ^ w44409;
	assign w24836 = w24752 ^ w24777;
	assign w24827 = w24828 ^ w24836;
	assign w24833 = w24834 ^ w24836;
	assign w24832 = w24835 & w24833;
	assign w24831 = w24832 ^ w24794;
	assign w24743 = w24832 ^ w24844;
	assign w24739 = w24743 ^ w24779;
	assign w24742 = w47245 ^ w24739;
	assign w24819 = w24741 ^ w24742;
	assign w24740 = w24832 ^ w24788;
	assign w24738 = w47247 ^ w24739;
	assign w24825 = w24836 & w24826;
	assign w24823 = w24825 ^ w24833;
	assign w24822 = w24831 & w24823;
	assign w24787 = w24822 ^ w24797;
	assign w24821 = w24787 ^ w24789;
	assign w24745 = w24822 ^ w24846;
	assign w24818 = w24787 ^ w24740;
	assign w24813 = w24827 & w47252;
	assign w24812 = w24818 & w24848;
	assign w24811 = w24821 & w24860;
	assign w24810 = w24831 & w24850;
	assign w24754 = w24810 ^ w24811;
	assign w24809 = w24819 & w24851;
	assign w24804 = w24827 & w24859;
	assign w24803 = w24818 & w24863;
	assign w24770 = w24812 ^ w24803;
	assign w24802 = w24821 & w24856;
	assign w24772 = w24810 ^ w24802;
	assign w24801 = w24831 & w24857;
	assign w24800 = w24819 & w24862;
	assign w44410 = w24811 ^ w24812;
	assign w44412 = w24825 ^ w24843;
	assign w24817 = w44412 ^ w24795;
	assign w24815 = w24817 & w24854;
	assign w44411 = w24813 ^ w24815;
	assign w24806 = w24817 & w24858;
	assign w24784 = w47251 ^ w44412;
	assign w24824 = w24784 ^ w24747;
	assign w24737 = w24784 ^ w24745;
	assign w24744 = w24774 ^ w24737;
	assign w24820 = w24741 ^ w24744;
	assign w24816 = w24737 ^ w24738;
	assign w24814 = w24824 & w24853;
	assign w24808 = w24816 & w24849;
	assign w24793 = w24808 ^ w44410;
	assign w24769 = w24808 ^ w24811;
	assign w24766 = ~w24769;
	assign w24765 = w24808 ^ w24809;
	assign w24759 = w24804 ^ w24793;
	assign w24756 = ~w24759;
	assign w24753 = w24809 ^ w24793;
	assign w24807 = w24820 & w24852;
	assign w24785 = w24803 ^ w24807;
	assign w24763 = ~w24785;
	assign w24762 = w24763 ^ w24801;
	assign w24758 = w24762 ^ w44411;
	assign w24761 = w24800 ^ w24758;
	assign w24805 = w24824 & w24855;
	assign w24799 = w24816 & w24864;
	assign w24798 = w24820 & w24861;
	assign w24764 = w24809 ^ w24798;
	assign w24760 = ~w24764;
	assign w24865 = w24760 ^ w24761;
	assign w43567 = w24799 ^ w24800;
	assign w24781 = w24805 ^ w43567;
	assign w24757 = w24781 ^ w24758;
	assign w49498 = w24756 ^ w24757;
	assign w24782 = w24806 ^ w24781;
	assign w49502 = w24782 ^ w24753;
	assign w24786 = w24814 ^ w24782;
	assign w24755 = w24813 ^ w24786;
	assign w49499 = w24754 ^ w24755;
	assign w24791 = w24815 ^ w24786;
	assign w24866 = w24791 ^ w24765;
	assign w49501 = ~w24866;
	assign w8457 = w49502 ^ w49514;
	assign w8213 = w8457 ^ w49498;
	assign w8533 = w8213 ^ w8214;
	assign w8471 = w49499 ^ w49512;
	assign w8256 = w8495 ^ w8457;
	assign w8442 = w8471 ^ w8462;
	assign w49500 = w44410 ^ w24791;
	assign w8251 = ~w49500;
	assign w8440 = w49513 ^ w8251;
	assign w24768 = w24772 ^ w43567;
	assign w24771 = w44411 ^ w24768;
	assign w24868 = w24770 ^ w24771;
	assign w24767 = w24763 ^ w24768;
	assign w24867 = w24766 ^ w24767;
	assign w45534 = ~w24734;
	assign w8244 = w8451 ^ w45534;
	assign w8520 = w8244 ^ w8245;
	assign w49339 = w8520 ^ w8493;
	assign w47099 = w49339 ^ w1844;
	assign w30759 = w47093 ^ w47099;
	assign w8515 = w45405 ^ w45534;
	assign w8383 = w8515 ^ w8493;
	assign w8267 = w8515 ^ w8452;
	assign w8392 = w8515 ^ w8453;
	assign w49322 = w45392 ^ w8267;
	assign w47116 = w49322 ^ w1827;
	assign w12452 = w47116 ^ w47110;
	assign w49330 = w45780 ^ w8392;
	assign w47108 = w49330 ^ w1835;
	assign w27594 = w47108 ^ w47102;
	assign w49314 = w45534 ^ w8444;
	assign w47124 = w49314 ^ w1819;
	assign w8321 = w49459 ^ w33709;
	assign w45538 = ~w24867;
	assign w8254 = w8463 ^ w45538;
	assign w45539 = ~w24868;
	assign w8211 = w8457 ^ w45539;
	assign w45540 = ~w24731;
	assign w8499 = w45390 ^ w45540;
	assign w8322 = w8499 ^ w49444;
	assign w8320 = ~w8322;
	assign w49319 = w8320 ^ w8321;
	assign w47119 = w49319 ^ w1824;
	assign w8304 = w45540 ^ w33710;
	assign w8302 = w8303 ^ w8304;
	assign w8395 = w8507 ^ w8499;
	assign w49327 = w45402 ^ w8395;
	assign w47111 = w49327 ^ w1832;
	assign w12532 = w47111 ^ w12452;
	assign w12446 = w47111 ^ w47109;
	assign w12529 = w12446 ^ w12452;
	assign w49320 = ~w8302;
	assign w47118 = w49320 ^ w1825;
	assign w17946 = w47124 ^ w47118;
	assign w17942 = w47120 ^ w47118;
	assign w17901 = w17942 ^ w47119;
	assign w18025 = w47124 ^ w17901;
	assign w18026 = w47119 ^ w17946;
	assign w18011 = w47124 & w18025;
	assign w8380 = w8504 ^ w45540;
	assign w49335 = w8380 ^ w8381;
	assign w47103 = w49335 ^ w1840;
	assign w27674 = w47103 ^ w27594;
	assign w27549 = w27590 ^ w47103;
	assign w27673 = w47108 ^ w27549;
	assign w27659 = w47108 & w27673;
	assign w45541 = ~w24733;
	assign w8373 = w45541 ^ w18167;
	assign w49340 = w8372 ^ w8373;
	assign w47098 = w49340 ^ w1845;
	assign w30686 = w47099 ^ w47098;
	assign w30757 = w47093 ^ w47098;
	assign w8384 = w8355 ^ w45541;
	assign w8514 = w45404 ^ w45541;
	assign w8390 = w8514 ^ w8492;
	assign w8367 = w8514 ^ w8491;
	assign w8389 = w8390 ^ w8391;
	assign w49316 = w49457 ^ w8367;
	assign w47122 = w49316 ^ w1821;
	assign w18030 = w47122 ^ w47120;
	assign w17916 = w47121 ^ w47122;
	assign w8382 = w8383 ^ w8384;
	assign w49315 = ~w8382;
	assign w47123 = w49315 ^ w1820;
	assign w17939 = w47123 ^ w47121;
	assign w17941 = w47122 ^ w17939;
	assign w18016 = w17946 ^ w17941;
	assign w17956 = w47123 ^ w47122;
	assign w18022 = w47123 ^ w18026;
	assign w18017 = w47118 ^ w17941;
	assign w18014 = w47119 ^ w17941;
	assign w18009 = w18026 & w18022;
	assign w45545 = ~w24865;
	assign w8424 = w24866 ^ w45545;
	assign w8480 = w45545 ^ w45535;
	assign w8438 = w8480 ^ w8468;
	assign w8414 = w8480 ^ w49509;
	assign w8366 = w8502 ^ w8499;
	assign w49344 = w45391 ^ w8366;
	assign w47094 = w49344 ^ w1849;
	assign w30676 = w47100 ^ w47094;
	assign w30753 = w30670 ^ w30676;
	assign w30751 = w30686 ^ w30753;
	assign w30756 = w47095 ^ w30676;
	assign w30752 = w47099 ^ w30756;
	assign w30739 = w30756 & w30752;
	assign w49331 = ~w8389;
	assign w47107 = w49331 ^ w1836;
	assign w27587 = w47107 ^ w47105;
	assign w27589 = w47106 ^ w27587;
	assign w27665 = w47102 ^ w27589;
	assign w27662 = w47103 ^ w27589;
	assign w27664 = w27594 ^ w27589;
	assign w27670 = w47107 ^ w27674;
	assign w27604 = w47107 ^ w47106;
	assign w27657 = w27674 & w27670;
	assign w45925 = ~w7971;
	assign w7873 = w45925 ^ w45417;
	assign w7871 = w7872 ^ w7873;
	assign w49154 = ~w7871;
	assign w47211 = w49154 ^ w1669;
	assign w12803 = w47205 ^ w47211;
	assign w12730 = w47211 ^ w47210;
	assign w12795 = w12730 ^ w12797;
	assign w7869 = w45925 ^ w49262;
	assign w49156 = w7868 ^ w7869;
	assign w47209 = w49156 ^ w1671;
	assign w12690 = w47209 ^ w47210;
	assign w12713 = w47211 ^ w47209;
	assign w12715 = w47210 ^ w12713;
	assign w12791 = w47206 ^ w12715;
	assign w12788 = w47207 ^ w12715;
	assign w12784 = w12803 & w12788;
	assign w12718 = w12784 ^ w12714;
	assign w12790 = w12720 ^ w12715;
	assign w12782 = w12797 & w12790;
	assign w7866 = w45925 ^ w49263;
	assign w49157 = w7865 ^ w7866;
	assign w47208 = w49157 ^ w1672;
	assign w12716 = w47208 ^ w47206;
	assign w12804 = w47210 ^ w47208;
	assign w12789 = w12714 ^ w12804;
	assign w12676 = w12716 ^ w12714;
	assign w12792 = w12713 ^ w12676;
	assign w12675 = w12716 ^ w47207;
	assign w12780 = w12804 & w12789;
	assign w12799 = w47212 ^ w12675;
	assign w12785 = w47212 & w12799;
	assign w12796 = w47211 ^ w12800;
	assign w12783 = w12800 & w12796;
	assign w12779 = w12801 & w12792;
	assign w43903 = w12779 ^ w12785;
	assign w12729 = w43903 ^ w12714;
	assign w43904 = w12779 ^ w12782;
	assign w12732 = w12780 ^ w43904;
	assign w12688 = w12783 ^ w12732;
	assign w12770 = w47211 ^ w12688;
	assign w12692 = w12718 ^ w43904;
	assign w12802 = w47208 ^ w47205;
	assign w12794 = w12713 ^ w12802;
	assign w12781 = w12802 & w12791;
	assign w12793 = w47212 ^ w12794;
	assign w12786 = w12795 & w12793;
	assign w12737 = w12780 ^ w12786;
	assign w12775 = w12737 ^ w12729;
	assign w12689 = w12780 ^ w12781;
	assign w12736 = w12689 ^ w12690;
	assign w12735 = w12736 ^ w12718;
	assign w12777 = w12783 ^ w12735;
	assign w12717 = w12781 ^ w12715;
	assign w12776 = w12692 ^ w12717;
	assign w12798 = w12802 ^ w12730;
	assign w12787 = w12794 & w12798;
	assign w12719 = w12787 ^ w12716;
	assign w12723 = w12719 ^ w12717;
	assign w12728 = w47205 ^ w12723;
	assign w12778 = w12737 ^ w12728;
	assign w12774 = w12778 & w12777;
	assign w12773 = w12774 ^ w12776;
	assign w12772 = w12775 & w12773;
	assign w12683 = w12772 ^ w12784;
	assign w12680 = w12772 ^ w12728;
	assign w12679 = w12683 ^ w12719;
	assign w12682 = w47205 ^ w12679;
	assign w12678 = w47207 ^ w12679;
	assign w12691 = w12723 ^ w43903;
	assign w12734 = w47207 ^ w12691;
	assign w12769 = w12774 ^ w12734;
	assign w12768 = w12769 & w12770;
	assign w12767 = w12768 ^ w12776;
	assign w12766 = w12774 ^ w12768;
	assign w12686 = w12768 ^ w12785;
	assign w12771 = w12772 ^ w12734;
	assign w12741 = w12771 & w12797;
	assign w12750 = w12771 & w12790;
	assign w12753 = w12767 & w47212;
	assign w12744 = w12767 & w12799;
	assign w12765 = w12776 & w12766;
	assign w12763 = w12765 ^ w12773;
	assign w12762 = w12771 & w12763;
	assign w12727 = w12762 ^ w12737;
	assign w12685 = w12762 ^ w12786;
	assign w12761 = w12727 ^ w12729;
	assign w12751 = w12761 & w12800;
	assign w12758 = w12727 ^ w12680;
	assign w12743 = w12758 & w12803;
	assign w12752 = w12758 & w12788;
	assign w12742 = w12761 & w12796;
	assign w12712 = w12750 ^ w12742;
	assign w43905 = w12751 ^ w12752;
	assign w12710 = w12752 ^ w12743;
	assign w12681 = w12686 ^ w12782;
	assign w12759 = w12681 ^ w12682;
	assign w12740 = w12759 & w12802;
	assign w12687 = w12768 ^ w12732;
	assign w43907 = w12765 ^ w12783;
	assign w12757 = w43907 ^ w12735;
	assign w12755 = w12757 & w12794;
	assign w43906 = w12753 ^ w12755;
	assign w12746 = w12757 & w12798;
	assign w12724 = w47211 ^ w43907;
	assign w12677 = w12724 ^ w12685;
	assign w12684 = w12714 ^ w12677;
	assign w12760 = w12681 ^ w12684;
	assign w12756 = w12677 ^ w12678;
	assign w12747 = w12760 & w12792;
	assign w12725 = w12743 ^ w12747;
	assign w12703 = ~w12725;
	assign w12739 = w12756 & w12804;
	assign w43532 = w12739 ^ w12740;
	assign w12708 = w12712 ^ w43532;
	assign w12711 = w43906 ^ w12708;
	assign w12808 = w12710 ^ w12711;
	assign w12707 = w12703 ^ w12708;
	assign w12738 = w12760 & w12801;
	assign w12702 = w12703 ^ w12741;
	assign w12698 = w12702 ^ w43906;
	assign w12764 = w12724 ^ w12687;
	assign w12754 = w12764 & w12793;
	assign w12701 = w12740 ^ w12698;
	assign w45250 = ~w12808;
	assign w8198 = w45397 ^ w45250;
	assign w8508 = w45539 ^ w45250;
	assign w8433 = w8508 ^ w8475;
	assign w49410 = w45250 ^ w8256;
	assign w8410 = w8508 ^ w8445;
	assign w49434 = w45397 ^ w8410;
	assign w47004 = w49434 ^ w1748;
	assign w47028 = w49410 ^ w1724;
	assign w12745 = w12764 & w12795;
	assign w12721 = w12745 ^ w43532;
	assign w12697 = w12721 ^ w12698;
	assign w12722 = w12746 ^ w12721;
	assign w12726 = w12754 ^ w12722;
	assign w12731 = w12755 ^ w12726;
	assign w49505 = w43905 ^ w12731;
	assign w8443 = w8457 ^ w49505;
	assign w8511 = w49500 ^ w49505;
	assign w49438 = w8517 ^ w8511;
	assign w47000 = w49438 ^ w1751;
	assign w49414 = w8442 ^ w8443;
	assign w47024 = w49414 ^ w1728;
	assign w12695 = w12753 ^ w12726;
	assign w8427 = w8511 ^ w8480;
	assign w49423 = w45394 ^ w8427;
	assign w47015 = w49423 ^ w1737;
	assign w12694 = w12750 ^ w12751;
	assign w49504 = w12694 ^ w12695;
	assign w8250 = w49504 ^ w8251;
	assign w8465 = w49504 ^ w49508;
	assign w49413 = w8533 ^ w8465;
	assign w47025 = w49413 ^ w1727;
	assign w8404 = w8465 ^ w8463;
	assign w8416 = w8511 ^ w8465;
	assign w12749 = w12759 & w12791;
	assign w12704 = w12749 ^ w12738;
	assign w12700 = ~w12704;
	assign w12805 = w12700 ^ w12701;
	assign w45255 = ~w12805;
	assign w8470 = w45255 ^ w45394;
	assign w8402 = w8470 ^ w8462;
	assign w8441 = ~w8470;
	assign w8415 = w45255 ^ w49505;
	assign w8423 = w8468 ^ w45255;
	assign w8422 = w8423 ^ w8424;
	assign w49424 = ~w8422;
	assign w47014 = w49424 ^ w1738;
	assign w8439 = w8441 ^ w45535;
	assign w49415 = w8439 ^ w8440;
	assign w49431 = w8414 ^ w8415;
	assign w47007 = w49431 ^ w1745;
	assign w49439 = w45545 ^ w8402;
	assign w47023 = w49415 ^ w1729;
	assign w46999 = w49439 ^ w1752;
	assign w12748 = w12756 & w12789;
	assign w12709 = w12748 ^ w12751;
	assign w12733 = w12748 ^ w43905;
	assign w12705 = w12748 ^ w12749;
	assign w12699 = w12744 ^ w12733;
	assign w12806 = w12731 ^ w12705;
	assign w12696 = ~w12699;
	assign w12706 = ~w12709;
	assign w12807 = w12706 ^ w12707;
	assign w49503 = w12696 ^ w12697;
	assign w8200 = w49504 ^ w49503;
	assign w8485 = w49498 ^ w49503;
	assign w8406 = w8485 ^ w8475;
	assign w49436 = w49507 ^ w8406;
	assign w47002 = w49436 ^ w45171;
	assign w17360 = w47002 ^ w47000;
	assign w8418 = w8485 ^ w49511;
	assign w8430 = w8485 ^ w8471;
	assign w8428 = ~w8430;
	assign w8255 = w45537 ^ w49503;
	assign w49412 = w8254 ^ w8255;
	assign w47026 = w49412 ^ w1726;
	assign w17494 = w47026 ^ w47024;
	assign w17380 = w47025 ^ w47026;
	assign w45256 = ~w12806;
	assign w8510 = w49501 ^ w45256;
	assign w8413 = w8510 ^ w8470;
	assign w8421 = w8510 ^ w8445;
	assign w49425 = w49502 ^ w8421;
	assign w8400 = w8510 ^ w45535;
	assign w49440 = w8400 ^ w8401;
	assign w46998 = w49440 ^ w1753;
	assign w17276 = w47004 ^ w46998;
	assign w17272 = w47000 ^ w46998;
	assign w17231 = w17272 ^ w46999;
	assign w17355 = w47004 ^ w17231;
	assign w49432 = w45536 ^ w8413;
	assign w8412 = w45395 ^ w45256;
	assign w17341 = w47004 & w17355;
	assign w47013 = w49425 ^ w1739;
	assign w12178 = w47015 ^ w47013;
	assign w49416 = w45256 ^ w8438;
	assign w47022 = w49416 ^ w1730;
	assign w17406 = w47024 ^ w47022;
	assign w17410 = w47028 ^ w47022;
	assign w17490 = w47023 ^ w17410;
	assign w17356 = w46999 ^ w17276;
	assign w45257 = ~w12807;
	assign w8212 = w45530 ^ w45257;
	assign w8500 = w45538 ^ w45257;
	assign w8431 = w8500 ^ w8463;
	assign w49420 = w49498 ^ w8431;
	assign w47018 = w49420 ^ w1734;
	assign w12265 = w47013 ^ w47018;
	assign w8534 = w8211 ^ w8212;
	assign w49411 = w8534 ^ w8475;
	assign w8419 = w45396 ^ w45257;
	assign w49428 = w8418 ^ w8419;
	assign w47010 = w49428 ^ w1742;
	assign w8409 = ~w8500;
	assign w8407 = w8409 ^ w8495;
	assign w47027 = w49411 ^ w1725;
	assign w17403 = w47027 ^ w47025;
	assign w17420 = w47027 ^ w47026;
	assign w17486 = w47027 ^ w17490;
	assign w17405 = w47026 ^ w17403;
	assign w17480 = w17410 ^ w17405;
	assign w17478 = w47023 ^ w17405;
	assign w17481 = w47022 ^ w17405;
	assign w17473 = w17490 & w17486;
	assign w17365 = w17406 ^ w47023;
	assign w17489 = w47028 ^ w17365;
	assign w17475 = w47028 & w17489;
	assign w12693 = w12749 ^ w12733;
	assign w49506 = w12722 ^ w12693;
	assign w8460 = w49506 ^ w49510;
	assign w8197 = w8460 ^ w45537;
	assign w8540 = w8197 ^ w8198;
	assign w8199 = w8460 ^ w49507;
	assign w8539 = w8199 ^ w8200;
	assign w8446 = w49502 ^ w49506;
	assign w49429 = w8539 ^ w8471;
	assign w47009 = w49429 ^ w1743;
	assign w24214 = w47009 ^ w47010;
	assign w8437 = w49506 ^ w24866;
	assign w8420 = w8508 ^ w8460;
	assign w49426 = w45530 ^ w8420;
	assign w8417 = w8460 ^ w49513;
	assign w49430 = w8416 ^ w8417;
	assign w47008 = w49430 ^ w1744;
	assign w24328 = w47010 ^ w47008;
	assign w47012 = w49426 ^ w1740;
	assign w8435 = w8495 ^ w8446;
	assign w8411 = w8446 ^ w49514;
	assign w49433 = w8411 ^ w8412;
	assign w47005 = w49433 ^ w1747;
	assign w24238 = w47007 ^ w47005;
	assign w24313 = w24238 ^ w24328;
	assign w24326 = w47008 ^ w47005;
	assign w24325 = w47005 ^ w47010;
	assign w24304 = w24328 & w24313;
	assign w8399 = w8468 ^ w8446;
	assign w49441 = w49510 ^ w8399;
	assign w49427 = w8540 ^ w8500;
	assign w47011 = w49427 ^ w1741;
	assign w24237 = w47011 ^ w47009;
	assign w24239 = w47010 ^ w24237;
	assign w24312 = w47007 ^ w24239;
	assign w24318 = w24237 ^ w24326;
	assign w24317 = w47012 ^ w24318;
	assign w24254 = w47011 ^ w47010;
	assign w24322 = w24326 ^ w24254;
	assign w24327 = w47005 ^ w47011;
	assign w24311 = w24318 & w24322;
	assign w24308 = w24327 & w24312;
	assign w24242 = w24308 ^ w24238;
	assign w49418 = w45539 ^ w8435;
	assign w47020 = w49418 ^ w1732;
	assign w12184 = w47020 ^ w47014;
	assign w12264 = w47015 ^ w12184;
	assign w12261 = w12178 ^ w12184;
	assign w46997 = w49441 ^ w1754;
	assign w17358 = w47000 ^ w46997;
	assign w17270 = w46999 ^ w46997;
	assign w17353 = w17270 ^ w17276;
	assign w17232 = w17272 ^ w17270;
	assign w17357 = w46997 ^ w47002;
	assign w17345 = w17270 ^ w17360;
	assign w17336 = w17360 & w17345;
	assign w47006 = w49432 ^ w1746;
	assign w24315 = w47006 ^ w24239;
	assign w24240 = w47008 ^ w47006;
	assign w24243 = w24311 ^ w24240;
	assign w24244 = w47012 ^ w47006;
	assign w24314 = w24244 ^ w24239;
	assign w24321 = w24238 ^ w24244;
	assign w24319 = w24254 ^ w24321;
	assign w24324 = w47007 ^ w24244;
	assign w24320 = w47011 ^ w24324;
	assign w24200 = w24240 ^ w24238;
	assign w24316 = w24237 ^ w24200;
	assign w24199 = w24240 ^ w47007;
	assign w24323 = w47012 ^ w24199;
	assign w24310 = w24319 & w24317;
	assign w24261 = w24304 ^ w24310;
	assign w24309 = w47012 & w24323;
	assign w24307 = w24324 & w24320;
	assign w24306 = w24321 & w24314;
	assign w24305 = w24326 & w24315;
	assign w24241 = w24305 ^ w24239;
	assign w24247 = w24243 ^ w24241;
	assign w24252 = w47005 ^ w24247;
	assign w24302 = w24261 ^ w24252;
	assign w24213 = w24304 ^ w24305;
	assign w24260 = w24213 ^ w24214;
	assign w24259 = w24260 ^ w24242;
	assign w24301 = w24307 ^ w24259;
	assign w24303 = w24325 & w24316;
	assign w24298 = w24302 & w24301;
	assign w44385 = w24303 ^ w24309;
	assign w24215 = w24247 ^ w44385;
	assign w24258 = w47007 ^ w24215;
	assign w24293 = w24298 ^ w24258;
	assign w24253 = w44385 ^ w24238;
	assign w24299 = w24261 ^ w24253;
	assign w44386 = w24303 ^ w24306;
	assign w24256 = w24304 ^ w44386;
	assign w24212 = w24307 ^ w24256;
	assign w24294 = w47011 ^ w24212;
	assign w24292 = w24293 & w24294;
	assign w24211 = w24292 ^ w24256;
	assign w24290 = w24298 ^ w24292;
	assign w24210 = w24292 ^ w24309;
	assign w24205 = w24210 ^ w24306;
	assign w24216 = w24242 ^ w44386;
	assign w24300 = w24216 ^ w24241;
	assign w24291 = w24292 ^ w24300;
	assign w24297 = w24298 ^ w24300;
	assign w24296 = w24299 & w24297;
	assign w24295 = w24296 ^ w24258;
	assign w24207 = w24296 ^ w24308;
	assign w24203 = w24207 ^ w24243;
	assign w24206 = w47005 ^ w24203;
	assign w24283 = w24205 ^ w24206;
	assign w24204 = w24296 ^ w24252;
	assign w24202 = w47007 ^ w24203;
	assign w24289 = w24300 & w24290;
	assign w24287 = w24289 ^ w24297;
	assign w24286 = w24295 & w24287;
	assign w24251 = w24286 ^ w24261;
	assign w24285 = w24251 ^ w24253;
	assign w24209 = w24286 ^ w24310;
	assign w24282 = w24251 ^ w24204;
	assign w24277 = w24291 & w47012;
	assign w24276 = w24282 & w24312;
	assign w24275 = w24285 & w24324;
	assign w24274 = w24295 & w24314;
	assign w24218 = w24274 ^ w24275;
	assign w24273 = w24283 & w24315;
	assign w24268 = w24291 & w24323;
	assign w24267 = w24282 & w24327;
	assign w24234 = w24276 ^ w24267;
	assign w24266 = w24285 & w24320;
	assign w24236 = w24274 ^ w24266;
	assign w24265 = w24295 & w24321;
	assign w24264 = w24283 & w24326;
	assign w44388 = w24275 ^ w24276;
	assign w44390 = w24289 ^ w24307;
	assign w24281 = w44390 ^ w24259;
	assign w24279 = w24281 & w24318;
	assign w44389 = w24277 ^ w24279;
	assign w24270 = w24281 & w24322;
	assign w24248 = w47011 ^ w44390;
	assign w24288 = w24248 ^ w24211;
	assign w24201 = w24248 ^ w24209;
	assign w24208 = w24238 ^ w24201;
	assign w24284 = w24205 ^ w24208;
	assign w24280 = w24201 ^ w24202;
	assign w24278 = w24288 & w24317;
	assign w24272 = w24280 & w24313;
	assign w24257 = w24272 ^ w44388;
	assign w24233 = w24272 ^ w24275;
	assign w24230 = ~w24233;
	assign w24229 = w24272 ^ w24273;
	assign w24223 = w24268 ^ w24257;
	assign w24220 = ~w24223;
	assign w24217 = w24273 ^ w24257;
	assign w24271 = w24284 & w24316;
	assign w24249 = w24267 ^ w24271;
	assign w24227 = ~w24249;
	assign w24226 = w24227 ^ w24265;
	assign w24222 = w24226 ^ w44389;
	assign w24225 = w24264 ^ w24222;
	assign w24269 = w24288 & w24319;
	assign w24263 = w24280 & w24328;
	assign w24262 = w24284 & w24325;
	assign w24228 = w24273 ^ w24262;
	assign w24224 = ~w24228;
	assign w24329 = w24224 ^ w24225;
	assign w44387 = w24263 ^ w24264;
	assign w24245 = w24269 ^ w44387;
	assign w24221 = w24245 ^ w24222;
	assign w49654 = w24220 ^ w24221;
	assign w24246 = w24270 ^ w24245;
	assign w49657 = w24246 ^ w24217;
	assign w24250 = w24278 ^ w24246;
	assign w24219 = w24277 ^ w24250;
	assign w49655 = w24218 ^ w24219;
	assign w24255 = w24279 ^ w24250;
	assign w24330 = w24255 ^ w24229;
	assign w8592 = ~w49654;
	assign w8591 = w49655 ^ w8592;
	assign w8770 = w45382 ^ w8592;
	assign w49656 = w44388 ^ w24255;
	assign w24232 = w24236 ^ w44387;
	assign w24235 = w44389 ^ w24232;
	assign w24332 = w24234 ^ w24235;
	assign w24231 = w24227 ^ w24232;
	assign w24331 = w24230 ^ w24231;
	assign w49653 = ~w24331;
	assign w8585 = w24331 ^ w45383;
	assign w45527 = ~w24329;
	assign w45528 = ~w24330;
	assign w45529 = ~w24332;
	assign w8589 = w45382 ^ w45529;
	assign w45926 = ~w7969;
	assign w7783 = w45926 ^ w49291;
	assign w49205 = w7782 ^ w7783;
	assign w47160 = w49205 ^ w1656;
	assign w30806 = w47160 ^ w47158;
	assign w30892 = w47160 ^ w47157;
	assign w30894 = w47162 ^ w47160;
	assign w30879 = w30804 ^ w30894;
	assign w30766 = w30806 ^ w30804;
	assign w30765 = w30806 ^ w47159;
	assign w30889 = w47164 ^ w30765;
	assign w30875 = w47164 & w30889;
	assign w30870 = w30894 & w30879;
	assign w7791 = w45926 ^ w45421;
	assign w49202 = w7790 ^ w7791;
	assign w47163 = w49202 ^ w1653;
	assign w30886 = w47163 ^ w30890;
	assign w30820 = w47163 ^ w47162;
	assign w30885 = w30820 ^ w30887;
	assign w30888 = w30892 ^ w30820;
	assign w30893 = w47157 ^ w47163;
	assign w30873 = w30890 & w30886;
	assign w7786 = w45926 ^ w49290;
	assign w49204 = w7785 ^ w7786;
	assign w47161 = w49204 ^ w1655;
	assign w30803 = w47163 ^ w47161;
	assign w30805 = w47162 ^ w30803;
	assign w30881 = w47158 ^ w30805;
	assign w30878 = w47159 ^ w30805;
	assign w30880 = w30810 ^ w30805;
	assign w30884 = w30803 ^ w30892;
	assign w30883 = w47164 ^ w30884;
	assign w30780 = w47161 ^ w47162;
	assign w30882 = w30803 ^ w30766;
	assign w30877 = w30884 & w30888;
	assign w30809 = w30877 ^ w30806;
	assign w30876 = w30885 & w30883;
	assign w30827 = w30870 ^ w30876;
	assign w30874 = w30893 & w30878;
	assign w30808 = w30874 ^ w30804;
	assign w30872 = w30887 & w30880;
	assign w30871 = w30892 & w30881;
	assign w30807 = w30871 ^ w30805;
	assign w30813 = w30809 ^ w30807;
	assign w30818 = w47157 ^ w30813;
	assign w30868 = w30827 ^ w30818;
	assign w30779 = w30870 ^ w30871;
	assign w30826 = w30779 ^ w30780;
	assign w30825 = w30826 ^ w30808;
	assign w30867 = w30873 ^ w30825;
	assign w30869 = w30891 & w30882;
	assign w30864 = w30868 & w30867;
	assign w44660 = w30869 ^ w30872;
	assign w30782 = w30808 ^ w44660;
	assign w30866 = w30782 ^ w30807;
	assign w30863 = w30864 ^ w30866;
	assign w30822 = w30870 ^ w44660;
	assign w30778 = w30873 ^ w30822;
	assign w30860 = w47163 ^ w30778;
	assign w44663 = w30869 ^ w30875;
	assign w30781 = w30813 ^ w44663;
	assign w30824 = w47159 ^ w30781;
	assign w30859 = w30864 ^ w30824;
	assign w30858 = w30859 & w30860;
	assign w30856 = w30864 ^ w30858;
	assign w30777 = w30858 ^ w30822;
	assign w30776 = w30858 ^ w30875;
	assign w30771 = w30776 ^ w30872;
	assign w30855 = w30866 & w30856;
	assign w30853 = w30855 ^ w30863;
	assign w44662 = w30855 ^ w30873;
	assign w30847 = w44662 ^ w30825;
	assign w30836 = w30847 & w30888;
	assign w30845 = w30847 & w30884;
	assign w30814 = w47163 ^ w44662;
	assign w30854 = w30814 ^ w30777;
	assign w30844 = w30854 & w30883;
	assign w30835 = w30854 & w30885;
	assign w30857 = w30858 ^ w30866;
	assign w30843 = w30857 & w47164;
	assign w30834 = w30857 & w30889;
	assign w30819 = w44663 ^ w30804;
	assign w30865 = w30827 ^ w30819;
	assign w30862 = w30865 & w30863;
	assign w30861 = w30862 ^ w30824;
	assign w30773 = w30862 ^ w30874;
	assign w30769 = w30773 ^ w30809;
	assign w30772 = w47157 ^ w30769;
	assign w30849 = w30771 ^ w30772;
	assign w30770 = w30862 ^ w30818;
	assign w30768 = w47159 ^ w30769;
	assign w30852 = w30861 & w30853;
	assign w30817 = w30852 ^ w30827;
	assign w30851 = w30817 ^ w30819;
	assign w30775 = w30852 ^ w30876;
	assign w30767 = w30814 ^ w30775;
	assign w30774 = w30804 ^ w30767;
	assign w30850 = w30771 ^ w30774;
	assign w30848 = w30817 ^ w30770;
	assign w30846 = w30767 ^ w30768;
	assign w30842 = w30848 & w30878;
	assign w30841 = w30851 & w30890;
	assign w30840 = w30861 & w30880;
	assign w30784 = w30840 ^ w30841;
	assign w30839 = w30849 & w30881;
	assign w30838 = w30846 & w30879;
	assign w30799 = w30838 ^ w30841;
	assign w30796 = ~w30799;
	assign w30795 = w30838 ^ w30839;
	assign w30837 = w30850 & w30882;
	assign w30833 = w30848 & w30893;
	assign w30815 = w30833 ^ w30837;
	assign w30800 = w30842 ^ w30833;
	assign w30793 = ~w30815;
	assign w30832 = w30851 & w30886;
	assign w30802 = w30840 ^ w30832;
	assign w30831 = w30861 & w30887;
	assign w30792 = w30793 ^ w30831;
	assign w30830 = w30849 & w30892;
	assign w30829 = w30846 & w30894;
	assign w30828 = w30850 & w30891;
	assign w30794 = w30839 ^ w30828;
	assign w30790 = ~w30794;
	assign w44661 = w30829 ^ w30830;
	assign w30811 = w30835 ^ w44661;
	assign w30812 = w30836 ^ w30811;
	assign w30816 = w30844 ^ w30812;
	assign w30785 = w30843 ^ w30816;
	assign w49495 = w30784 ^ w30785;
	assign w8487 = w49491 ^ w49495;
	assign w8290 = w8281 ^ w8487;
	assign w8232 = w8235 ^ w49495;
	assign w8525 = w8232 ^ w8233;
	assign w8260 = w8262 ^ w8487;
	assign w49389 = w8290 ^ w8291;
	assign w49397 = w8525 ^ w8498;
	assign w47041 = w49397 ^ w1774;
	assign w47049 = w49389 ^ w1766;
	assign w30821 = w30845 ^ w30816;
	assign w30896 = w30821 ^ w30795;
	assign w30798 = w30802 ^ w44661;
	assign w30797 = w30793 ^ w30798;
	assign w30897 = w30796 ^ w30797;
	assign w44664 = w30841 ^ w30842;
	assign w49496 = w44664 ^ w30821;
	assign w8478 = w49492 ^ w49496;
	assign w8288 = w8265 ^ w8478;
	assign w49390 = w8288 ^ w8289;
	assign w47048 = w49390 ^ w1767;
	assign w8259 = w8483 ^ w8478;
	assign w49407 = w45633 ^ w8259;
	assign w47031 = w49407 ^ w1784;
	assign w8236 = w8235 ^ w49496;
	assign w8524 = w8236 ^ w8237;
	assign w49398 = w8524 ^ w8490;
	assign w47040 = w49398 ^ w1775;
	assign w30823 = w30838 ^ w44664;
	assign w30789 = w30834 ^ w30823;
	assign w30786 = ~w30789;
	assign w30783 = w30839 ^ w30823;
	assign w49497 = w30812 ^ w30783;
	assign w8447 = w49493 ^ w49497;
	assign w8455 = w49482 ^ w49497;
	assign w8228 = w8455 ^ w49495;
	assign w8224 = ~w8455;
	assign w8272 = w45891 ^ w49497;
	assign w49401 = w8272 ^ w8273;
	assign w47037 = w49401 ^ w1778;
	assign w17626 = w47040 ^ w47037;
	assign w8271 = w8513 ^ w8447;
	assign w49402 = w45628 ^ w8271;
	assign w47036 = w49402 ^ w1779;
	assign w8285 = w8476 ^ w8447;
	assign w49393 = w49482 ^ w8285;
	assign w47045 = w49393 ^ w1770;
	assign w12400 = w47048 ^ w47045;
	assign w44665 = w30843 ^ w30845;
	assign w30801 = w44665 ^ w30798;
	assign w30898 = w30800 ^ w30801;
	assign w30788 = w30792 ^ w44665;
	assign w30791 = w30830 ^ w30788;
	assign w30895 = w30790 ^ w30791;
	assign w30787 = w30811 ^ w30788;
	assign w49494 = w30786 ^ w30787;
	assign w8279 = w8281 ^ w49494;
	assign w8497 = w49490 ^ w49494;
	assign w8292 = w8512 ^ w8497;
	assign w49388 = w49479 ^ w8292;
	assign w49396 = w8279 ^ w8280;
	assign w8263 = w8265 ^ w8497;
	assign w47050 = w49388 ^ w1765;
	assign w47042 = w49396 ^ w1773;
	assign w17628 = w47042 ^ w47040;
	assign w17514 = w47041 ^ w47042;
	assign w17625 = w47037 ^ w47042;
	assign w12288 = w47049 ^ w47050;
	assign w12402 = w47050 ^ w47048;
	assign w12399 = w47045 ^ w47050;
	assign w8225 = w8224 ^ w49494;
	assign w8528 = w8225 ^ w8226;
	assign w49381 = w8528 ^ w8487;
	assign w47057 = w49381 ^ w1758;
	assign w8310 = ~w8497;
	assign w8527 = w8228 ^ w8229;
	assign w49382 = w8527 ^ w8478;
	assign w47056 = w49382 ^ w1759;
	assign w45706 = ~w30897;
	assign w8308 = w8310 ^ w45706;
	assign w49380 = w8308 ^ w8309;
	assign w8230 = w8454 ^ w45706;
	assign w8526 = w8230 ^ w8231;
	assign w49395 = w8526 ^ w8512;
	assign w47043 = w49395 ^ w1772;
	assign w17537 = w47043 ^ w47041;
	assign w17539 = w47042 ^ w17537;
	assign w17627 = w47037 ^ w47043;
	assign w17618 = w17537 ^ w17626;
	assign w17554 = w47043 ^ w47042;
	assign w47058 = w49380 ^ w1757;
	assign w27544 = w47058 ^ w47056;
	assign w27430 = w47057 ^ w47058;
	assign w8501 = w45627 ^ w45706;
	assign w8266 = w8505 ^ w8501;
	assign w49404 = w49490 ^ w8266;
	assign w8294 = w8513 ^ w8501;
	assign w8293 = w8294 ^ w8295;
	assign w49387 = ~w8293;
	assign w47051 = w49387 ^ w1764;
	assign w12328 = w47051 ^ w47050;
	assign w12401 = w47045 ^ w47051;
	assign w12311 = w47051 ^ w47049;
	assign w12392 = w12311 ^ w12400;
	assign w12396 = w12400 ^ w12328;
	assign w12313 = w47050 ^ w12311;
	assign w12385 = w12392 & w12396;
	assign w47034 = w49404 ^ w1781;
	assign w17622 = w17626 ^ w17554;
	assign w17611 = w17618 & w17622;
	assign w45707 = ~w30898;
	assign w8509 = w45628 ^ w45707;
	assign w8270 = w8512 ^ w8509;
	assign w8268 = ~w8270;
	assign w8296 = w8509 ^ w8450;
	assign w49386 = w45624 ^ w8296;
	assign w8222 = w8224 ^ w45707;
	assign w8529 = w8222 ^ w8223;
	assign w49379 = w8529 ^ w8501;
	assign w47059 = w49379 ^ w1756;
	assign w27453 = w47059 ^ w47057;
	assign w27455 = w47058 ^ w27453;
	assign w27470 = w47059 ^ w47058;
	assign w47052 = w49386 ^ w1763;
	assign w12391 = w47052 ^ w12392;
	assign w49394 = w45707 ^ w8282;
	assign w47044 = w49394 ^ w1771;
	assign w17617 = w47044 ^ w17618;
	assign w8311 = w8509 ^ w8455;
	assign w49378 = w45254 ^ w8311;
	assign w47060 = w49378 ^ w1755;
	assign w45712 = ~w30895;
	assign w8472 = w45633 ^ w45712;
	assign w8287 = w8490 ^ w8472;
	assign w49391 = w45629 ^ w8287;
	assign w47047 = w49391 ^ w1768;
	assign w8307 = w8472 ^ w49496;
	assign w8305 = ~w8307;
	assign w49383 = w8305 ^ w8306;
	assign w47055 = w49383 ^ w1760;
	assign w27528 = w47055 ^ w27455;
	assign w12312 = w47047 ^ w47045;
	assign w12387 = w12312 ^ w12402;
	assign w12378 = w12402 & w12387;
	assign w12386 = w47047 ^ w12313;
	assign w12382 = w12401 & w12386;
	assign w12316 = w12382 ^ w12312;
	assign w8258 = w8476 ^ w8472;
	assign w49408 = w45626 ^ w8258;
	assign w47030 = w49408 ^ w1785;
	assign w24378 = w47036 ^ w47030;
	assign w24458 = w47031 ^ w24378;
	assign w8277 = w8483 ^ w45712;
	assign w49399 = w8277 ^ w8278;
	assign w47039 = w49399 ^ w1776;
	assign w17612 = w47039 ^ w17539;
	assign w17538 = w47039 ^ w47037;
	assign w17613 = w17538 ^ w17628;
	assign w17608 = w17627 & w17612;
	assign w17542 = w17608 ^ w17538;
	assign w17604 = w17628 & w17613;
	assign w45713 = ~w30896;
	assign w8297 = w8447 ^ w45713;
	assign w49385 = w8297 ^ w8298;
	assign w8461 = w45626 ^ w45713;
	assign w8286 = w8483 ^ w8461;
	assign w49392 = w45622 ^ w8286;
	assign w47053 = w49385 ^ w1762;
	assign w27454 = w47055 ^ w47053;
	assign w27529 = w27454 ^ w27544;
	assign w27542 = w47056 ^ w47053;
	assign w27538 = w27542 ^ w27470;
	assign w27534 = w27453 ^ w27542;
	assign w27533 = w47060 ^ w27534;
	assign w27543 = w47053 ^ w47059;
	assign w27541 = w47053 ^ w47058;
	assign w27527 = w27534 & w27538;
	assign w27524 = w27543 & w27528;
	assign w27458 = w27524 ^ w27454;
	assign w27520 = w27544 & w27529;
	assign w47046 = w49392 ^ w1769;
	assign w12318 = w47052 ^ w47046;
	assign w12388 = w12318 ^ w12313;
	assign w12398 = w47047 ^ w12318;
	assign w12395 = w12312 ^ w12318;
	assign w12380 = w12395 & w12388;
	assign w12394 = w47051 ^ w12398;
	assign w12393 = w12328 ^ w12395;
	assign w12384 = w12393 & w12391;
	assign w12381 = w12398 & w12394;
	assign w12335 = w12378 ^ w12384;
	assign w12389 = w47046 ^ w12313;
	assign w12379 = w12400 & w12389;
	assign w12315 = w12379 ^ w12313;
	assign w12287 = w12378 ^ w12379;
	assign w12334 = w12287 ^ w12288;
	assign w12333 = w12334 ^ w12316;
	assign w12375 = w12381 ^ w12333;
	assign w12314 = w47048 ^ w47046;
	assign w12317 = w12385 ^ w12314;
	assign w12274 = w12314 ^ w12312;
	assign w12321 = w12317 ^ w12315;
	assign w12326 = w47045 ^ w12321;
	assign w12376 = w12335 ^ w12326;
	assign w12390 = w12311 ^ w12274;
	assign w12273 = w12314 ^ w47047;
	assign w12397 = w47052 ^ w12273;
	assign w12383 = w47052 & w12397;
	assign w12377 = w12399 & w12390;
	assign w12372 = w12376 & w12375;
	assign w8276 = w8476 ^ w45713;
	assign w8274 = ~w8276;
	assign w49400 = w8274 ^ w8275;
	assign w47038 = w49400 ^ w1777;
	assign w17615 = w47038 ^ w17539;
	assign w17540 = w47040 ^ w47038;
	assign w17543 = w17611 ^ w17540;
	assign w17500 = w17540 ^ w17538;
	assign w17616 = w17537 ^ w17500;
	assign w17499 = w17540 ^ w47039;
	assign w17623 = w47044 ^ w17499;
	assign w17609 = w47044 & w17623;
	assign w17544 = w47044 ^ w47038;
	assign w17624 = w47039 ^ w17544;
	assign w17620 = w47043 ^ w17624;
	assign w17614 = w17544 ^ w17539;
	assign w17621 = w17538 ^ w17544;
	assign w17619 = w17554 ^ w17621;
	assign w17610 = w17619 & w17617;
	assign w17561 = w17604 ^ w17610;
	assign w17607 = w17624 & w17620;
	assign w17606 = w17621 & w17614;
	assign w17605 = w17626 & w17615;
	assign w17513 = w17604 ^ w17605;
	assign w17560 = w17513 ^ w17514;
	assign w17559 = w17560 ^ w17542;
	assign w17541 = w17605 ^ w17539;
	assign w17547 = w17543 ^ w17541;
	assign w17552 = w47037 ^ w17547;
	assign w17602 = w17561 ^ w17552;
	assign w17601 = w17607 ^ w17559;
	assign w17603 = w17625 & w17616;
	assign w17598 = w17602 & w17601;
	assign w8257 = w8461 ^ w8450;
	assign w49409 = w49493 ^ w8257;
	assign w47029 = w49409 ^ w1786;
	assign w24459 = w47029 ^ w47034;
	assign w24372 = w47031 ^ w47029;
	assign w8300 = w8461 ^ w45712;
	assign w43886 = w12377 ^ w12383;
	assign w12327 = w43886 ^ w12312;
	assign w12373 = w12335 ^ w12327;
	assign w12289 = w12321 ^ w43886;
	assign w12332 = w47047 ^ w12289;
	assign w12367 = w12372 ^ w12332;
	assign w43887 = w12377 ^ w12380;
	assign w12330 = w12378 ^ w43887;
	assign w12286 = w12381 ^ w12330;
	assign w12368 = w47051 ^ w12286;
	assign w12366 = w12367 & w12368;
	assign w12364 = w12372 ^ w12366;
	assign w12285 = w12366 ^ w12330;
	assign w12284 = w12366 ^ w12383;
	assign w12279 = w12284 ^ w12380;
	assign w12290 = w12316 ^ w43887;
	assign w12374 = w12290 ^ w12315;
	assign w12371 = w12372 ^ w12374;
	assign w12370 = w12373 & w12371;
	assign w12369 = w12370 ^ w12332;
	assign w12339 = w12369 & w12395;
	assign w12278 = w12370 ^ w12326;
	assign w12281 = w12370 ^ w12382;
	assign w12277 = w12281 ^ w12317;
	assign w12276 = w47047 ^ w12277;
	assign w12280 = w47045 ^ w12277;
	assign w12357 = w12279 ^ w12280;
	assign w12338 = w12357 & w12400;
	assign w12363 = w12374 & w12364;
	assign w12361 = w12363 ^ w12371;
	assign w12360 = w12369 & w12361;
	assign w12325 = w12360 ^ w12335;
	assign w12359 = w12325 ^ w12327;
	assign w12340 = w12359 & w12394;
	assign w12356 = w12325 ^ w12278;
	assign w12350 = w12356 & w12386;
	assign w12349 = w12359 & w12398;
	assign w12283 = w12360 ^ w12384;
	assign w12341 = w12356 & w12401;
	assign w12308 = w12350 ^ w12341;
	assign w12365 = w12366 ^ w12374;
	assign w12351 = w12365 & w47052;
	assign w12342 = w12365 & w12397;
	assign w43888 = w12349 ^ w12350;
	assign w43890 = w12363 ^ w12381;
	assign w12322 = w47051 ^ w43890;
	assign w12362 = w12322 ^ w12285;
	assign w12343 = w12362 & w12393;
	assign w12275 = w12322 ^ w12283;
	assign w12354 = w12275 ^ w12276;
	assign w12346 = w12354 & w12387;
	assign w12337 = w12354 & w12402;
	assign w12307 = w12346 ^ w12349;
	assign w12304 = ~w12307;
	assign w12282 = w12312 ^ w12275;
	assign w12358 = w12279 ^ w12282;
	assign w12336 = w12358 & w12399;
	assign w12345 = w12358 & w12390;
	assign w12323 = w12341 ^ w12345;
	assign w12301 = ~w12323;
	assign w12300 = w12301 ^ w12339;
	assign w43531 = w12337 ^ w12338;
	assign w12319 = w12343 ^ w43531;
	assign w12352 = w12362 & w12391;
	assign w12331 = w12346 ^ w43888;
	assign w12297 = w12342 ^ w12331;
	assign w12294 = ~w12297;
	assign w12355 = w43890 ^ w12333;
	assign w12344 = w12355 & w12396;
	assign w12320 = w12344 ^ w12319;
	assign w12324 = w12352 ^ w12320;
	assign w12353 = w12355 & w12392;
	assign w12329 = w12353 ^ w12324;
	assign w49649 = w43888 ^ w12329;
	assign w8851 = w49645 ^ w49649;
	assign w12293 = w12351 ^ w12324;
	assign w8725 = w49656 ^ w49649;
	assign w43889 = w12351 ^ w12353;
	assign w12296 = w12300 ^ w43889;
	assign w12299 = w12338 ^ w12296;
	assign w12295 = w12319 ^ w12296;
	assign w49647 = w12294 ^ w12295;
	assign w8835 = w49647 ^ w49654;
	assign w8587 = w49643 ^ w49647;
	assign w8718 = ~w8835;
	assign w8716 = w8718 ^ w49643;
	assign w44103 = w17603 ^ w17609;
	assign w17515 = w17547 ^ w44103;
	assign w17558 = w47039 ^ w17515;
	assign w17593 = w17598 ^ w17558;
	assign w17553 = w44103 ^ w17538;
	assign w17599 = w17561 ^ w17553;
	assign w44104 = w17603 ^ w17606;
	assign w17556 = w17604 ^ w44104;
	assign w17512 = w17607 ^ w17556;
	assign w17594 = w47043 ^ w17512;
	assign w17592 = w17593 & w17594;
	assign w17590 = w17598 ^ w17592;
	assign w17510 = w17592 ^ w17609;
	assign w17505 = w17510 ^ w17606;
	assign w17511 = w17592 ^ w17556;
	assign w17516 = w17542 ^ w44104;
	assign w17600 = w17516 ^ w17541;
	assign w17597 = w17598 ^ w17600;
	assign w17591 = w17592 ^ w17600;
	assign w17577 = w17591 & w47044;
	assign w17596 = w17599 & w17597;
	assign w17504 = w17596 ^ w17552;
	assign w17595 = w17596 ^ w17558;
	assign w17507 = w17596 ^ w17608;
	assign w17503 = w17507 ^ w17543;
	assign w17502 = w47039 ^ w17503;
	assign w17506 = w47037 ^ w17503;
	assign w17583 = w17505 ^ w17506;
	assign w17573 = w17583 & w17615;
	assign w17574 = w17595 & w17614;
	assign w17565 = w17595 & w17621;
	assign w17568 = w17591 & w17623;
	assign w8299 = w8300 ^ w8301;
	assign w49384 = ~w8299;
	assign w47054 = w49384 ^ w1761;
	assign w27531 = w47054 ^ w27455;
	assign w27456 = w47056 ^ w47054;
	assign w27459 = w27527 ^ w27456;
	assign w27460 = w47060 ^ w47054;
	assign w27530 = w27460 ^ w27455;
	assign w27537 = w27454 ^ w27460;
	assign w27535 = w27470 ^ w27537;
	assign w27540 = w47055 ^ w27460;
	assign w27536 = w47059 ^ w27540;
	assign w27416 = w27456 ^ w27454;
	assign w27532 = w27453 ^ w27416;
	assign w27415 = w27456 ^ w47055;
	assign w27539 = w47060 ^ w27415;
	assign w27526 = w27535 & w27533;
	assign w27477 = w27520 ^ w27526;
	assign w27525 = w47060 & w27539;
	assign w27523 = w27540 & w27536;
	assign w27522 = w27537 & w27530;
	assign w27521 = w27542 & w27531;
	assign w27457 = w27521 ^ w27455;
	assign w27463 = w27459 ^ w27457;
	assign w27468 = w47053 ^ w27463;
	assign w27518 = w27477 ^ w27468;
	assign w27429 = w27520 ^ w27521;
	assign w27476 = w27429 ^ w27430;
	assign w27475 = w27476 ^ w27458;
	assign w27517 = w27523 ^ w27475;
	assign w27519 = w27541 & w27532;
	assign w27514 = w27518 & w27517;
	assign w44518 = w27519 ^ w27525;
	assign w27469 = w44518 ^ w27454;
	assign w27515 = w27477 ^ w27469;
	assign w27431 = w27463 ^ w44518;
	assign w27474 = w47055 ^ w27431;
	assign w27509 = w27514 ^ w27474;
	assign w44519 = w27519 ^ w27522;
	assign w27472 = w27520 ^ w44519;
	assign w27428 = w27523 ^ w27472;
	assign w27510 = w47059 ^ w27428;
	assign w27508 = w27509 & w27510;
	assign w27427 = w27508 ^ w27472;
	assign w27426 = w27508 ^ w27525;
	assign w27421 = w27426 ^ w27522;
	assign w27506 = w27514 ^ w27508;
	assign w27432 = w27458 ^ w44519;
	assign w27516 = w27432 ^ w27457;
	assign w27507 = w27508 ^ w27516;
	assign w27513 = w27514 ^ w27516;
	assign w27512 = w27515 & w27513;
	assign w27511 = w27512 ^ w27474;
	assign w27423 = w27512 ^ w27524;
	assign w27419 = w27423 ^ w27459;
	assign w27422 = w47053 ^ w27419;
	assign w27499 = w27421 ^ w27422;
	assign w27420 = w27512 ^ w27468;
	assign w27418 = w47055 ^ w27419;
	assign w27505 = w27516 & w27506;
	assign w27503 = w27505 ^ w27513;
	assign w27502 = w27511 & w27503;
	assign w27467 = w27502 ^ w27477;
	assign w27501 = w27467 ^ w27469;
	assign w27425 = w27502 ^ w27526;
	assign w27498 = w27467 ^ w27420;
	assign w27493 = w27507 & w47060;
	assign w27492 = w27498 & w27528;
	assign w27491 = w27501 & w27540;
	assign w27490 = w27511 & w27530;
	assign w27434 = w27490 ^ w27491;
	assign w27489 = w27499 & w27531;
	assign w27484 = w27507 & w27539;
	assign w27483 = w27498 & w27543;
	assign w27450 = w27492 ^ w27483;
	assign w27482 = w27501 & w27536;
	assign w27452 = w27490 ^ w27482;
	assign w27481 = w27511 & w27537;
	assign w27480 = w27499 & w27542;
	assign w44520 = w27491 ^ w27492;
	assign w44522 = w27505 ^ w27523;
	assign w27464 = w47059 ^ w44522;
	assign w27504 = w27464 ^ w27427;
	assign w27485 = w27504 & w27535;
	assign w27494 = w27504 & w27533;
	assign w27417 = w27464 ^ w27425;
	assign w27424 = w27454 ^ w27417;
	assign w27500 = w27421 ^ w27424;
	assign w27487 = w27500 & w27532;
	assign w27465 = w27483 ^ w27487;
	assign w27443 = ~w27465;
	assign w27442 = w27443 ^ w27481;
	assign w27496 = w27417 ^ w27418;
	assign w27479 = w27496 & w27544;
	assign w27478 = w27500 & w27541;
	assign w27444 = w27489 ^ w27478;
	assign w27440 = ~w27444;
	assign w43577 = w27479 ^ w27480;
	assign w27461 = w27485 ^ w43577;
	assign w27448 = w27452 ^ w43577;
	assign w27447 = w27443 ^ w27448;
	assign w27488 = w27496 & w27529;
	assign w27449 = w27488 ^ w27491;
	assign w27446 = ~w27449;
	assign w27547 = w27446 ^ w27447;
	assign w27445 = w27488 ^ w27489;
	assign w27473 = w27488 ^ w44520;
	assign w27433 = w27489 ^ w27473;
	assign w27439 = w27484 ^ w27473;
	assign w27436 = ~w27439;
	assign w27497 = w44522 ^ w27475;
	assign w27495 = w27497 & w27534;
	assign w27486 = w27497 & w27538;
	assign w27462 = w27486 ^ w27461;
	assign w27466 = w27494 ^ w27462;
	assign w27471 = w27495 ^ w27466;
	assign w49665 = w44520 ^ w27471;
	assign w27546 = w27471 ^ w27445;
	assign w27435 = w27493 ^ w27466;
	assign w49664 = w27434 ^ w27435;
	assign w49666 = w27462 ^ w27433;
	assign w8802 = w49666 ^ w49679;
	assign w8549 = ~w8802;
	assign w8550 = w8549 ^ w49676;
	assign w8547 = w8549 ^ w45698;
	assign w8553 = w8802 ^ w49677;
	assign w44521 = w27493 ^ w27495;
	assign w27451 = w44521 ^ w27448;
	assign w27548 = w27450 ^ w27451;
	assign w27438 = w27442 ^ w44521;
	assign w27441 = w27480 ^ w27438;
	assign w27545 = w27440 ^ w27441;
	assign w27437 = w27461 ^ w27438;
	assign w49663 = w27436 ^ w27437;
	assign w17589 = w17600 & w17590;
	assign w17587 = w17589 ^ w17597;
	assign w17586 = w17595 & w17587;
	assign w17509 = w17586 ^ w17610;
	assign w17551 = w17586 ^ w17561;
	assign w17582 = w17551 ^ w17504;
	assign w17576 = w17582 & w17612;
	assign w17585 = w17551 ^ w17553;
	assign w17566 = w17585 & w17620;
	assign w17536 = w17574 ^ w17566;
	assign w44108 = w17589 ^ w17607;
	assign w17548 = w47043 ^ w44108;
	assign w17588 = w17548 ^ w17511;
	assign w17578 = w17588 & w17617;
	assign w17501 = w17548 ^ w17509;
	assign w17508 = w17538 ^ w17501;
	assign w17584 = w17505 ^ w17508;
	assign w17562 = w17584 & w17625;
	assign w17528 = w17573 ^ w17562;
	assign w17524 = ~w17528;
	assign w17580 = w17501 ^ w17502;
	assign w17563 = w17580 & w17628;
	assign w17572 = w17580 & w17613;
	assign w17529 = w17572 ^ w17573;
	assign w17581 = w44108 ^ w17559;
	assign w17579 = w17581 & w17618;
	assign w17570 = w17581 & w17622;
	assign w44107 = w17577 ^ w17579;
	assign w12348 = w12369 & w12388;
	assign w12310 = w12348 ^ w12340;
	assign w12292 = w12348 ^ w12349;
	assign w49648 = w12292 ^ w12293;
	assign w8860 = w49644 ^ w49648;
	assign w12306 = w12310 ^ w43531;
	assign w12305 = w12301 ^ w12306;
	assign w12405 = w12304 ^ w12305;
	assign w8583 = w49655 ^ w49648;
	assign w8729 = w8860 ^ w8718;
	assign w8742 = ~w8860;
	assign w12309 = w43889 ^ w12306;
	assign w12406 = w12308 ^ w12309;
	assign w12347 = w12357 & w12389;
	assign w12303 = w12346 ^ w12347;
	assign w12404 = w12329 ^ w12303;
	assign w49651 = ~w12404;
	assign w8846 = w45389 ^ w49651;
	assign w12291 = w12347 ^ w12331;
	assign w49652 = w12320 ^ w12291;
	assign w8796 = w49646 ^ w49652;
	assign w8797 = w49652 ^ w49657;
	assign w8586 = w8796 ^ w49644;
	assign w8865 = w8586 ^ w8587;
	assign w8721 = w45528 ^ w12404;
	assign w8731 = ~w8797;
	assign w12302 = w12347 ^ w12336;
	assign w12298 = ~w12302;
	assign w12403 = w12298 ^ w12299;
	assign w49650 = ~w12403;
	assign w8848 = w45388 ^ w49650;
	assign w8723 = w45527 ^ w12403;
	assign w17569 = w17588 & w17619;
	assign w45247 = ~w12405;
	assign w8837 = w45247 ^ w49653;
	assign w8735 = w8731 ^ w45247;
	assign w45248 = ~w12406;
	assign w8836 = w45248 ^ w45529;
	assign w24455 = w24372 ^ w24378;
	assign w45614 = ~w27546;
	assign w8811 = w45614 ^ w45704;
	assign w8684 = w49666 ^ w45614;
	assign w45615 = ~w27547;
	assign w45616 = ~w27548;
	assign w45621 = ~w27545;
	assign w8703 = w45703 ^ w45621;
	assign w17575 = w17585 & w17624;
	assign w17518 = w17574 ^ w17575;
	assign w17533 = w17572 ^ w17575;
	assign w17530 = ~w17533;
	assign w44106 = w17575 ^ w17576;
	assign w17557 = w17572 ^ w44106;
	assign w17523 = w17568 ^ w17557;
	assign w17517 = w17573 ^ w17557;
	assign w17520 = ~w17523;
	assign w17571 = w17584 & w17616;
	assign w17567 = w17582 & w17627;
	assign w17549 = w17567 ^ w17571;
	assign w17527 = ~w17549;
	assign w17526 = w17527 ^ w17565;
	assign w17534 = w17576 ^ w17567;
	assign w17522 = w17526 ^ w44107;
	assign w17564 = w17583 & w17626;
	assign w17525 = w17564 ^ w17522;
	assign w17629 = w17524 ^ w17525;
	assign w44105 = w17563 ^ w17564;
	assign w17545 = w17569 ^ w44105;
	assign w17546 = w17570 ^ w17545;
	assign w49711 = w17546 ^ w17517;
	assign w17550 = w17578 ^ w17546;
	assign w17555 = w17579 ^ w17550;
	assign w49710 = w44106 ^ w17555;
	assign w17630 = w17555 ^ w17529;
	assign w17519 = w17577 ^ w17550;
	assign w49709 = w17518 ^ w17519;
	assign w8597 = w49710 ^ w49709;
	assign w17532 = w17536 ^ w44105;
	assign w17535 = w44107 ^ w17532;
	assign w17632 = w17534 ^ w17535;
	assign w17531 = w17527 ^ w17532;
	assign w17631 = w17530 ^ w17531;
	assign w17521 = w17545 ^ w17522;
	assign w49708 = w17520 ^ w17521;
	assign w45374 = ~w17631;
	assign w45375 = ~w17632;
	assign w45380 = ~w17629;
	assign w45381 = ~w17630;
	assign w8745 = w45381 ^ w45380;
	assign w45927 = ~w8449;
	assign w8344 = w45927 ^ w49464;
	assign w49358 = w8343 ^ w8344;
	assign w47080 = w49358 ^ w1799;
	assign w33486 = w47080 ^ w47078;
	assign w33572 = w47080 ^ w47077;
	assign w33574 = w47082 ^ w47080;
	assign w33559 = w33484 ^ w33574;
	assign w33446 = w33486 ^ w33484;
	assign w33445 = w33486 ^ w47079;
	assign w33569 = w47084 ^ w33445;
	assign w33555 = w47084 & w33569;
	assign w33550 = w33574 & w33559;
	assign w8351 = w45927 ^ w45400;
	assign w8349 = w8350 ^ w8351;
	assign w49355 = ~w8349;
	assign w47083 = w49355 ^ w1796;
	assign w33566 = w47083 ^ w33570;
	assign w33500 = w47083 ^ w47082;
	assign w33565 = w33500 ^ w33567;
	assign w33568 = w33572 ^ w33500;
	assign w33573 = w47077 ^ w47083;
	assign w33553 = w33570 & w33566;
	assign w8347 = w45927 ^ w49463;
	assign w49357 = w8346 ^ w8347;
	assign w47081 = w49357 ^ w1798;
	assign w33483 = w47083 ^ w47081;
	assign w33485 = w47082 ^ w33483;
	assign w33561 = w47078 ^ w33485;
	assign w33558 = w47079 ^ w33485;
	assign w33560 = w33490 ^ w33485;
	assign w33564 = w33483 ^ w33572;
	assign w33563 = w47084 ^ w33564;
	assign w33460 = w47081 ^ w47082;
	assign w33562 = w33483 ^ w33446;
	assign w33557 = w33564 & w33568;
	assign w33489 = w33557 ^ w33486;
	assign w33556 = w33565 & w33563;
	assign w33507 = w33550 ^ w33556;
	assign w33554 = w33573 & w33558;
	assign w33488 = w33554 ^ w33484;
	assign w33552 = w33567 & w33560;
	assign w33551 = w33572 & w33561;
	assign w33487 = w33551 ^ w33485;
	assign w33493 = w33489 ^ w33487;
	assign w33498 = w47077 ^ w33493;
	assign w33548 = w33507 ^ w33498;
	assign w33459 = w33550 ^ w33551;
	assign w33506 = w33459 ^ w33460;
	assign w33505 = w33506 ^ w33488;
	assign w33547 = w33553 ^ w33505;
	assign w33549 = w33571 & w33562;
	assign w33544 = w33548 & w33547;
	assign w44771 = w33549 ^ w33552;
	assign w33462 = w33488 ^ w44771;
	assign w33546 = w33462 ^ w33487;
	assign w33543 = w33544 ^ w33546;
	assign w33502 = w33550 ^ w44771;
	assign w33458 = w33553 ^ w33502;
	assign w33540 = w47083 ^ w33458;
	assign w44774 = w33549 ^ w33555;
	assign w33461 = w33493 ^ w44774;
	assign w33504 = w47079 ^ w33461;
	assign w33539 = w33544 ^ w33504;
	assign w33538 = w33539 & w33540;
	assign w33536 = w33544 ^ w33538;
	assign w33457 = w33538 ^ w33502;
	assign w33456 = w33538 ^ w33555;
	assign w33451 = w33456 ^ w33552;
	assign w33535 = w33546 & w33536;
	assign w33533 = w33535 ^ w33543;
	assign w44773 = w33535 ^ w33553;
	assign w33527 = w44773 ^ w33505;
	assign w33516 = w33527 & w33568;
	assign w33525 = w33527 & w33564;
	assign w33494 = w47083 ^ w44773;
	assign w33534 = w33494 ^ w33457;
	assign w33524 = w33534 & w33563;
	assign w33515 = w33534 & w33565;
	assign w33537 = w33538 ^ w33546;
	assign w33523 = w33537 & w47084;
	assign w33514 = w33537 & w33569;
	assign w33499 = w44774 ^ w33484;
	assign w33545 = w33507 ^ w33499;
	assign w33542 = w33545 & w33543;
	assign w33541 = w33542 ^ w33504;
	assign w33453 = w33542 ^ w33554;
	assign w33449 = w33453 ^ w33489;
	assign w33452 = w47077 ^ w33449;
	assign w33529 = w33451 ^ w33452;
	assign w33450 = w33542 ^ w33498;
	assign w33448 = w47079 ^ w33449;
	assign w33532 = w33541 & w33533;
	assign w33497 = w33532 ^ w33507;
	assign w33531 = w33497 ^ w33499;
	assign w33455 = w33532 ^ w33556;
	assign w33447 = w33494 ^ w33455;
	assign w33454 = w33484 ^ w33447;
	assign w33530 = w33451 ^ w33454;
	assign w33528 = w33497 ^ w33450;
	assign w33526 = w33447 ^ w33448;
	assign w33522 = w33528 & w33558;
	assign w33521 = w33531 & w33570;
	assign w33520 = w33541 & w33560;
	assign w33464 = w33520 ^ w33521;
	assign w33519 = w33529 & w33561;
	assign w33518 = w33526 & w33559;
	assign w33479 = w33518 ^ w33521;
	assign w33476 = ~w33479;
	assign w33475 = w33518 ^ w33519;
	assign w33517 = w33530 & w33562;
	assign w33513 = w33528 & w33573;
	assign w33495 = w33513 ^ w33517;
	assign w33480 = w33522 ^ w33513;
	assign w33473 = ~w33495;
	assign w33512 = w33531 & w33566;
	assign w33482 = w33520 ^ w33512;
	assign w33511 = w33541 & w33567;
	assign w33472 = w33473 ^ w33511;
	assign w33510 = w33529 & w33572;
	assign w33509 = w33526 & w33574;
	assign w33508 = w33530 & w33571;
	assign w33474 = w33519 ^ w33508;
	assign w33470 = ~w33474;
	assign w44772 = w33509 ^ w33510;
	assign w33491 = w33515 ^ w44772;
	assign w33492 = w33516 ^ w33491;
	assign w33496 = w33524 ^ w33492;
	assign w33465 = w33523 ^ w33496;
	assign w49705 = w33464 ^ w33465;
	assign w8809 = w49705 ^ w49709;
	assign w33501 = w33525 ^ w33496;
	assign w33576 = w33501 ^ w33475;
	assign w33478 = w33482 ^ w44772;
	assign w33477 = w33473 ^ w33478;
	assign w33577 = w33476 ^ w33477;
	assign w44775 = w33521 ^ w33522;
	assign w49706 = w44775 ^ w33501;
	assign w33503 = w33518 ^ w44775;
	assign w33469 = w33514 ^ w33503;
	assign w33466 = ~w33469;
	assign w33463 = w33519 ^ w33503;
	assign w49707 = w33492 ^ w33463;
	assign w8804 = w49707 ^ w49711;
	assign w8543 = w8804 ^ w49708;
	assign w44776 = w33523 ^ w33525;
	assign w33481 = w44776 ^ w33478;
	assign w33578 = w33480 ^ w33481;
	assign w33468 = w33472 ^ w44776;
	assign w33471 = w33510 ^ w33468;
	assign w33575 = w33470 ^ w33471;
	assign w33467 = w33491 ^ w33468;
	assign w49704 = w33466 ^ w33467;
	assign w8544 = w49705 ^ w49704;
	assign w8883 = w8543 ^ w8544;
	assign w45774 = ~w33576;
	assign w8756 = w45381 ^ w45774;
	assign w45775 = ~w33577;
	assign w8763 = w45374 ^ w45775;
	assign w45776 = ~w33578;
	assign w8542 = w45375 ^ w45776;
	assign w45781 = ~w33575;
	assign w8814 = w45781 ^ w45380;
	assign w8785 = ~w8814;
	assign w8759 = w45781 ^ w49706;
	assign w45928 = ~w8447;
	assign w8269 = w45928 ^ w45627;
	assign w49403 = w8268 ^ w8269;
	assign w47035 = w49403 ^ w1780;
	assign w24388 = w47035 ^ w47034;
	assign w24454 = w47035 ^ w24458;
	assign w24461 = w47029 ^ w47035;
	assign w24441 = w24458 & w24454;
	assign w24453 = w24388 ^ w24455;
	assign w8264 = w45928 ^ w49491;
	assign w49405 = w8263 ^ w8264;
	assign w47033 = w49405 ^ w1782;
	assign w24348 = w47033 ^ w47034;
	assign w24371 = w47035 ^ w47033;
	assign w24373 = w47034 ^ w24371;
	assign w24449 = w47030 ^ w24373;
	assign w24446 = w47031 ^ w24373;
	assign w24448 = w24378 ^ w24373;
	assign w24442 = w24461 & w24446;
	assign w24376 = w24442 ^ w24372;
	assign w24440 = w24455 & w24448;
	assign w8261 = w45928 ^ w49492;
	assign w49406 = w8260 ^ w8261;
	assign w47032 = w49406 ^ w1783;
	assign w24374 = w47032 ^ w47030;
	assign w24333 = w24374 ^ w47031;
	assign w24457 = w47036 ^ w24333;
	assign w24334 = w24374 ^ w24372;
	assign w24450 = w24371 ^ w24334;
	assign w24437 = w24459 & w24450;
	assign w24460 = w47032 ^ w47029;
	assign w24456 = w24460 ^ w24388;
	assign w24439 = w24460 & w24449;
	assign w24375 = w24439 ^ w24373;
	assign w24443 = w47036 & w24457;
	assign w44391 = w24437 ^ w24443;
	assign w24387 = w44391 ^ w24372;
	assign w24462 = w47034 ^ w47032;
	assign w24447 = w24372 ^ w24462;
	assign w24438 = w24462 & w24447;
	assign w24347 = w24438 ^ w24439;
	assign w24394 = w24347 ^ w24348;
	assign w24393 = w24394 ^ w24376;
	assign w24435 = w24441 ^ w24393;
	assign w44392 = w24437 ^ w24440;
	assign w24350 = w24376 ^ w44392;
	assign w24434 = w24350 ^ w24375;
	assign w24390 = w24438 ^ w44392;
	assign w24346 = w24441 ^ w24390;
	assign w24428 = w47035 ^ w24346;
	assign w24452 = w24371 ^ w24460;
	assign w24451 = w47036 ^ w24452;
	assign w24444 = w24453 & w24451;
	assign w24445 = w24452 & w24456;
	assign w24377 = w24445 ^ w24374;
	assign w24381 = w24377 ^ w24375;
	assign w24349 = w24381 ^ w44391;
	assign w24392 = w47031 ^ w24349;
	assign w24395 = w24438 ^ w24444;
	assign w24433 = w24395 ^ w24387;
	assign w24386 = w47029 ^ w24381;
	assign w24436 = w24395 ^ w24386;
	assign w24432 = w24436 & w24435;
	assign w24427 = w24432 ^ w24392;
	assign w24431 = w24432 ^ w24434;
	assign w24426 = w24427 & w24428;
	assign w24344 = w24426 ^ w24443;
	assign w24345 = w24426 ^ w24390;
	assign w24339 = w24344 ^ w24440;
	assign w24425 = w24426 ^ w24434;
	assign w24402 = w24425 & w24457;
	assign w24411 = w24425 & w47036;
	assign w24430 = w24433 & w24431;
	assign w24341 = w24430 ^ w24442;
	assign w24338 = w24430 ^ w24386;
	assign w24337 = w24341 ^ w24377;
	assign w24340 = w47029 ^ w24337;
	assign w24417 = w24339 ^ w24340;
	assign w24398 = w24417 & w24460;
	assign w24336 = w47031 ^ w24337;
	assign w24407 = w24417 & w24449;
	assign w24424 = w24432 ^ w24426;
	assign w24423 = w24434 & w24424;
	assign w24421 = w24423 ^ w24431;
	assign w24429 = w24430 ^ w24392;
	assign w24399 = w24429 & w24455;
	assign w24420 = w24429 & w24421;
	assign w24385 = w24420 ^ w24395;
	assign w24408 = w24429 & w24448;
	assign w24416 = w24385 ^ w24338;
	assign w24401 = w24416 & w24461;
	assign w24410 = w24416 & w24446;
	assign w24368 = w24410 ^ w24401;
	assign w24419 = w24385 ^ w24387;
	assign w24400 = w24419 & w24454;
	assign w24370 = w24408 ^ w24400;
	assign w24409 = w24419 & w24458;
	assign w24352 = w24408 ^ w24409;
	assign w24343 = w24420 ^ w24444;
	assign w44393 = w24409 ^ w24410;
	assign w44395 = w24423 ^ w24441;
	assign w24382 = w47035 ^ w44395;
	assign w24335 = w24382 ^ w24343;
	assign w24342 = w24372 ^ w24335;
	assign w24418 = w24339 ^ w24342;
	assign w24396 = w24418 & w24459;
	assign w24414 = w24335 ^ w24336;
	assign w24397 = w24414 & w24462;
	assign w24406 = w24414 & w24447;
	assign w24363 = w24406 ^ w24407;
	assign w24367 = w24406 ^ w24409;
	assign w24364 = ~w24367;
	assign w24405 = w24418 & w24450;
	assign w24383 = w24401 ^ w24405;
	assign w24361 = ~w24383;
	assign w24360 = w24361 ^ w24399;
	assign w24362 = w24407 ^ w24396;
	assign w24358 = ~w24362;
	assign w43566 = w24397 ^ w24398;
	assign w24366 = w24370 ^ w43566;
	assign w24365 = w24361 ^ w24366;
	assign w24465 = w24364 ^ w24365;
	assign w24422 = w24382 ^ w24345;
	assign w24403 = w24422 & w24453;
	assign w24379 = w24403 ^ w43566;
	assign w24391 = w24406 ^ w44393;
	assign w24351 = w24407 ^ w24391;
	assign w24357 = w24402 ^ w24391;
	assign w24354 = ~w24357;
	assign w24412 = w24422 & w24451;
	assign w24415 = w44395 ^ w24393;
	assign w24404 = w24415 & w24456;
	assign w24413 = w24415 & w24452;
	assign w24380 = w24404 ^ w24379;
	assign w49698 = w24380 ^ w24351;
	assign w8791 = w49694 ^ w49698;
	assign w24384 = w24412 ^ w24380;
	assign w24389 = w24413 ^ w24384;
	assign w24464 = w24389 ^ w24363;
	assign w24353 = w24411 ^ w24384;
	assign w49696 = w24352 ^ w24353;
	assign w8831 = w49692 ^ w49696;
	assign w44394 = w24411 ^ w24413;
	assign w24369 = w44394 ^ w24366;
	assign w24466 = w24368 ^ w24369;
	assign w24356 = w24360 ^ w44394;
	assign w24359 = w24398 ^ w24356;
	assign w24463 = w24358 ^ w24359;
	assign w24355 = w24379 ^ w24356;
	assign w49697 = w44393 ^ w24389;
	assign w8822 = w49693 ^ w49697;
	assign w45526 = ~w24466;
	assign w8853 = w45379 ^ w45526;
	assign w45531 = ~w24463;
	assign w8816 = w45384 ^ w45531;
	assign w8651 = w8816 ^ w49697;
	assign w8649 = ~w8651;
	assign w45532 = ~w24464;
	assign w8805 = w45385 ^ w45532;
	assign w8644 = w8805 ^ w45531;
	assign w8641 = w8791 ^ w45532;
	assign w45533 = ~w24465;
	assign w8845 = w45378 ^ w45533;
	assign w49695 = w24354 ^ w24355;
	assign w8841 = w49691 ^ w49695;
	assign w8654 = ~w8841;
	assign w8652 = w8654 ^ w45533;
	assign w45929 = ~w8446;
	assign w8434 = w45929 ^ w45538;
	assign w8429 = w45929 ^ w49508;
	assign w8249 = w45929 ^ w49499;
	assign w8518 = w8249 ^ w8250;
	assign w49422 = w8518 ^ w8462;
	assign w47016 = w49422 ^ w1736;
	assign w12268 = w47018 ^ w47016;
	assign w12266 = w47016 ^ w47013;
	assign w12253 = w12178 ^ w12268;
	assign w12244 = w12268 & w12253;
	assign w49421 = w8428 ^ w8429;
	assign w8432 = w8433 ^ w8434;
	assign w49419 = ~w8432;
	assign w47019 = w49419 ^ w1733;
	assign w12267 = w47013 ^ w47019;
	assign w12260 = w47019 ^ w12264;
	assign w12247 = w12264 & w12260;
	assign w12194 = w47019 ^ w47018;
	assign w12259 = w12194 ^ w12261;
	assign w12262 = w12266 ^ w12194;
	assign w12180 = w47016 ^ w47014;
	assign w12139 = w12180 ^ w47015;
	assign w12263 = w47020 ^ w12139;
	assign w12140 = w12180 ^ w12178;
	assign w12249 = w47020 & w12263;
	assign w47017 = w49421 ^ w1735;
	assign w12154 = w47017 ^ w47018;
	assign w12177 = w47019 ^ w47017;
	assign w12258 = w12177 ^ w12266;
	assign w12257 = w47020 ^ w12258;
	assign w12256 = w12177 ^ w12140;
	assign w12243 = w12265 & w12256;
	assign w12251 = w12258 & w12262;
	assign w12183 = w12251 ^ w12180;
	assign w12250 = w12259 & w12257;
	assign w12179 = w47018 ^ w12177;
	assign w12255 = w47014 ^ w12179;
	assign w12254 = w12184 ^ w12179;
	assign w12246 = w12261 & w12254;
	assign w12201 = w12244 ^ w12250;
	assign w43880 = w12243 ^ w12249;
	assign w12193 = w43880 ^ w12178;
	assign w12239 = w12201 ^ w12193;
	assign w12245 = w12266 & w12255;
	assign w12153 = w12244 ^ w12245;
	assign w12200 = w12153 ^ w12154;
	assign w43881 = w12243 ^ w12246;
	assign w12196 = w12244 ^ w43881;
	assign w12152 = w12247 ^ w12196;
	assign w12234 = w47019 ^ w12152;
	assign w12181 = w12245 ^ w12179;
	assign w12187 = w12183 ^ w12181;
	assign w12192 = w47013 ^ w12187;
	assign w12155 = w12187 ^ w43880;
	assign w12198 = w47015 ^ w12155;
	assign w12242 = w12201 ^ w12192;
	assign w12252 = w47015 ^ w12179;
	assign w12248 = w12267 & w12252;
	assign w12182 = w12248 ^ w12178;
	assign w12156 = w12182 ^ w43881;
	assign w12240 = w12156 ^ w12181;
	assign w12199 = w12200 ^ w12182;
	assign w12241 = w12247 ^ w12199;
	assign w12238 = w12242 & w12241;
	assign w12233 = w12238 ^ w12198;
	assign w12232 = w12233 & w12234;
	assign w12231 = w12232 ^ w12240;
	assign w12237 = w12238 ^ w12240;
	assign w12151 = w12232 ^ w12196;
	assign w12217 = w12231 & w47020;
	assign w12236 = w12239 & w12237;
	assign w12147 = w12236 ^ w12248;
	assign w12143 = w12147 ^ w12183;
	assign w12146 = w47013 ^ w12143;
	assign w12142 = w47015 ^ w12143;
	assign w12150 = w12232 ^ w12249;
	assign w12145 = w12150 ^ w12246;
	assign w12223 = w12145 ^ w12146;
	assign w12213 = w12223 & w12255;
	assign w12230 = w12238 ^ w12232;
	assign w12229 = w12240 & w12230;
	assign w12227 = w12229 ^ w12237;
	assign w43885 = w12229 ^ w12247;
	assign w12221 = w43885 ^ w12199;
	assign w12219 = w12221 & w12258;
	assign w43884 = w12217 ^ w12219;
	assign w12188 = w47019 ^ w43885;
	assign w12228 = w12188 ^ w12151;
	assign w12218 = w12228 & w12257;
	assign w12144 = w12236 ^ w12192;
	assign w12210 = w12221 & w12262;
	assign w12209 = w12228 & w12259;
	assign w12208 = w12231 & w12263;
	assign w12204 = w12223 & w12266;
	assign w12235 = w12236 ^ w12198;
	assign w12226 = w12235 & w12227;
	assign w12214 = w12235 & w12254;
	assign w12149 = w12226 ^ w12250;
	assign w12141 = w12188 ^ w12149;
	assign w12148 = w12178 ^ w12141;
	assign w12220 = w12141 ^ w12142;
	assign w12224 = w12145 ^ w12148;
	assign w12211 = w12224 & w12256;
	assign w12212 = w12220 & w12253;
	assign w12169 = w12212 ^ w12213;
	assign w12205 = w12235 & w12261;
	assign w12203 = w12220 & w12268;
	assign w43882 = w12203 ^ w12204;
	assign w12185 = w12209 ^ w43882;
	assign w12186 = w12210 ^ w12185;
	assign w12190 = w12218 ^ w12186;
	assign w12159 = w12217 ^ w12190;
	assign w12195 = w12219 ^ w12190;
	assign w12270 = w12195 ^ w12169;
	assign w45242 = ~w12270;
	assign w12191 = w12226 ^ w12201;
	assign w12222 = w12191 ^ w12144;
	assign w12216 = w12222 & w12252;
	assign w12225 = w12191 ^ w12193;
	assign w12215 = w12225 & w12264;
	assign w12158 = w12214 ^ w12215;
	assign w49669 = w12158 ^ w12159;
	assign w8825 = w49664 ^ w49669;
	assign w8689 = ~w8825;
	assign w12173 = w12212 ^ w12215;
	assign w12170 = ~w12173;
	assign w12207 = w12222 & w12267;
	assign w12174 = w12216 ^ w12207;
	assign w12189 = w12207 ^ w12211;
	assign w43883 = w12215 ^ w12216;
	assign w12197 = w12212 ^ w43883;
	assign w12163 = w12208 ^ w12197;
	assign w12160 = ~w12163;
	assign w49670 = w43883 ^ w12195;
	assign w8554 = w49670 ^ w49664;
	assign w8879 = w8553 ^ w8554;
	assign w8821 = w49665 ^ w49670;
	assign w8663 = ~w8821;
	assign w12167 = ~w12189;
	assign w12166 = w12167 ^ w12205;
	assign w12162 = w12166 ^ w43884;
	assign w12161 = w12185 ^ w12162;
	assign w49668 = w12160 ^ w12161;
	assign w8828 = w49663 ^ w49668;
	assign w12165 = w12204 ^ w12162;
	assign w8681 = ~w8828;
	assign w8679 = w8681 ^ w49676;
	assign w8707 = w49668 ^ w45615;
	assign w12157 = w12213 ^ w12197;
	assign w49671 = w12186 ^ w12157;
	assign w8793 = w49666 ^ w49671;
	assign w8656 = w8793 ^ w45704;
	assign w8552 = ~w49669;
	assign w8551 = w8552 ^ w49663;
	assign w8880 = w8550 ^ w8551;
	assign w12206 = w12225 & w12260;
	assign w12176 = w12214 ^ w12206;
	assign w12172 = w12176 ^ w43882;
	assign w12175 = w43884 ^ w12172;
	assign w12272 = w12174 ^ w12175;
	assign w12171 = w12167 ^ w12172;
	assign w12271 = w12170 ^ w12171;
	assign w8548 = w12271 ^ w45616;
	assign w8881 = w8547 ^ w8548;
	assign w49667 = ~w12271;
	assign w8832 = w45615 ^ w49667;
	assign w45243 = ~w12272;
	assign w8833 = w45616 ^ w45243;
	assign w12202 = w12224 & w12265;
	assign w12168 = w12213 ^ w12202;
	assign w12164 = ~w12168;
	assign w12269 = w12164 ^ w12165;
	assign w45249 = ~w12269;
	assign w8675 = w45242 ^ w45249;
	assign w8705 = w45249 ^ w49665;
	assign w8817 = w45621 ^ w45249;
	assign w8685 = w8817 ^ w8811;
	assign w8678 = w8817 ^ w45703;
	assign w8676 = ~w8678;
	assign w45930 = ~w8445;
	assign w8408 = w45930 ^ w45396;
	assign w49435 = w8407 ^ w8408;
	assign w47003 = w49435 ^ w1749;
	assign w17359 = w46997 ^ w47003;
	assign w17286 = w47003 ^ w47002;
	assign w8436 = w45930 ^ w45536;
	assign w49417 = w8436 ^ w8437;
	assign w17351 = w17286 ^ w17353;
	assign w17354 = w17358 ^ w17286;
	assign w8405 = w45930 ^ w49499;
	assign w8403 = w8404 ^ w8405;
	assign w49437 = ~w8403;
	assign w17352 = w47003 ^ w17356;
	assign w17339 = w17356 & w17352;
	assign w47021 = w49417 ^ w1731;
	assign w17492 = w47024 ^ w47021;
	assign w17471 = w17492 & w17481;
	assign w17407 = w17471 ^ w17405;
	assign w17491 = w47021 ^ w47026;
	assign w17488 = w17492 ^ w17420;
	assign w17484 = w17403 ^ w17492;
	assign w17483 = w47028 ^ w17484;
	assign w17477 = w17484 & w17488;
	assign w17409 = w17477 ^ w17406;
	assign w17404 = w47023 ^ w47021;
	assign w17479 = w17404 ^ w17494;
	assign w17470 = w17494 & w17479;
	assign w17366 = w17406 ^ w17404;
	assign w17379 = w17470 ^ w17471;
	assign w17426 = w17379 ^ w17380;
	assign w17487 = w17404 ^ w17410;
	assign w17485 = w17420 ^ w17487;
	assign w17476 = w17485 & w17483;
	assign w17472 = w17487 & w17480;
	assign w17427 = w17470 ^ w17476;
	assign w17413 = w17409 ^ w17407;
	assign w17418 = w47021 ^ w17413;
	assign w17468 = w17427 ^ w17418;
	assign w47001 = w49437 ^ w1750;
	assign w17269 = w47003 ^ w47001;
	assign w17350 = w17269 ^ w17358;
	assign w17348 = w17269 ^ w17232;
	assign w17335 = w17357 & w17348;
	assign w17343 = w17350 & w17354;
	assign w17275 = w17343 ^ w17272;
	assign w17246 = w47001 ^ w47002;
	assign w17271 = w47002 ^ w17269;
	assign w17347 = w46998 ^ w17271;
	assign w17346 = w17276 ^ w17271;
	assign w17338 = w17353 & w17346;
	assign w17344 = w46999 ^ w17271;
	assign w17340 = w17359 & w17344;
	assign w17274 = w17340 ^ w17270;
	assign w17337 = w17358 & w17347;
	assign w17273 = w17337 ^ w17271;
	assign w17245 = w17336 ^ w17337;
	assign w17292 = w17245 ^ w17246;
	assign w17291 = w17292 ^ w17274;
	assign w17333 = w17339 ^ w17291;
	assign w17349 = w47004 ^ w17350;
	assign w17342 = w17351 & w17349;
	assign w17293 = w17336 ^ w17342;
	assign w44092 = w17335 ^ w17338;
	assign w17288 = w17336 ^ w44092;
	assign w17244 = w17339 ^ w17288;
	assign w17326 = w47003 ^ w17244;
	assign w44095 = w17335 ^ w17341;
	assign w17285 = w44095 ^ w17270;
	assign w17331 = w17293 ^ w17285;
	assign w17279 = w17275 ^ w17273;
	assign w17247 = w17279 ^ w44095;
	assign w17290 = w46999 ^ w17247;
	assign w17284 = w46997 ^ w17279;
	assign w17334 = w17293 ^ w17284;
	assign w17330 = w17334 & w17333;
	assign w17325 = w17330 ^ w17290;
	assign w17324 = w17325 & w17326;
	assign w17243 = w17324 ^ w17288;
	assign w17322 = w17330 ^ w17324;
	assign w17242 = w17324 ^ w17341;
	assign w17237 = w17242 ^ w17338;
	assign w17482 = w17403 ^ w17366;
	assign w17469 = w17491 & w17482;
	assign w44098 = w17469 ^ w17475;
	assign w17419 = w44098 ^ w17404;
	assign w17465 = w17427 ^ w17419;
	assign w17381 = w17413 ^ w44098;
	assign w17424 = w47023 ^ w17381;
	assign w44099 = w17469 ^ w17472;
	assign w17422 = w17470 ^ w44099;
	assign w17378 = w17473 ^ w17422;
	assign w17460 = w47027 ^ w17378;
	assign w17248 = w17274 ^ w44092;
	assign w17332 = w17248 ^ w17273;
	assign w17329 = w17330 ^ w17332;
	assign w17328 = w17331 & w17329;
	assign w17236 = w17328 ^ w17284;
	assign w17327 = w17328 ^ w17290;
	assign w17306 = w17327 & w17346;
	assign w17297 = w17327 & w17353;
	assign w17323 = w17324 ^ w17332;
	assign w17300 = w17323 & w17355;
	assign w17239 = w17328 ^ w17340;
	assign w17235 = w17239 ^ w17275;
	assign w17234 = w46999 ^ w17235;
	assign w17238 = w46997 ^ w17235;
	assign w17315 = w17237 ^ w17238;
	assign w17296 = w17315 & w17358;
	assign w17309 = w17323 & w47004;
	assign w17305 = w17315 & w17347;
	assign w17321 = w17332 & w17322;
	assign w17319 = w17321 ^ w17329;
	assign w17318 = w17327 & w17319;
	assign w17283 = w17318 ^ w17293;
	assign w17314 = w17283 ^ w17236;
	assign w17308 = w17314 & w17344;
	assign w17299 = w17314 & w17359;
	assign w17266 = w17308 ^ w17299;
	assign w17317 = w17283 ^ w17285;
	assign w17298 = w17317 & w17352;
	assign w17307 = w17317 & w17356;
	assign w17250 = w17306 ^ w17307;
	assign w17268 = w17306 ^ w17298;
	assign w44094 = w17321 ^ w17339;
	assign w17280 = w47003 ^ w44094;
	assign w17320 = w17280 ^ w17243;
	assign w17310 = w17320 & w17349;
	assign w17301 = w17320 & w17351;
	assign w44096 = w17307 ^ w17308;
	assign w17313 = w44094 ^ w17291;
	assign w17302 = w17313 & w17354;
	assign w17311 = w17313 & w17350;
	assign w44097 = w17309 ^ w17311;
	assign w17241 = w17318 ^ w17342;
	assign w17233 = w17280 ^ w17241;
	assign w17240 = w17270 ^ w17233;
	assign w17316 = w17237 ^ w17240;
	assign w17303 = w17316 & w17348;
	assign w17312 = w17233 ^ w17234;
	assign w17281 = w17299 ^ w17303;
	assign w17259 = ~w17281;
	assign w17258 = w17259 ^ w17297;
	assign w17254 = w17258 ^ w44097;
	assign w17257 = w17296 ^ w17254;
	assign w17304 = w17312 & w17345;
	assign w17261 = w17304 ^ w17305;
	assign w17289 = w17304 ^ w44096;
	assign w17265 = w17304 ^ w17307;
	assign w17262 = ~w17265;
	assign w17255 = w17300 ^ w17289;
	assign w17252 = ~w17255;
	assign w17294 = w17316 & w17357;
	assign w17260 = w17305 ^ w17294;
	assign w17256 = ~w17260;
	assign w17361 = w17256 ^ w17257;
	assign w17249 = w17305 ^ w17289;
	assign w17295 = w17312 & w17360;
	assign w44093 = w17295 ^ w17296;
	assign w45372 = ~w17361;
	assign w8783 = w8785 ^ w45372;
	assign w17277 = w17301 ^ w44093;
	assign w17253 = w17277 ^ w17254;
	assign w49712 = w17252 ^ w17253;
	assign w8807 = w49708 ^ w49712;
	assign w17278 = w17302 ^ w17277;
	assign w17282 = w17310 ^ w17278;
	assign w49715 = w17278 ^ w17249;
	assign w17251 = w17309 ^ w17282;
	assign w49713 = w17250 ^ w17251;
	assign w8558 = w49713 ^ w49712;
	assign w8748 = w8809 ^ w8807;
	assign w17287 = w17311 ^ w17282;
	assign w17362 = w17287 ^ w17261;
	assign w49714 = w44096 ^ w17287;
	assign w8806 = w49710 ^ w49714;
	assign w8746 = w8814 ^ w8806;
	assign w8761 = w8804 ^ w49714;
	assign w8789 = w49711 ^ w49715;
	assign w8596 = w8789 ^ w49713;
	assign w8861 = w8596 ^ w8597;
	assign w45373 = ~w17362;
	assign w8812 = w45381 ^ w45373;
	assign w8767 = w8812 ^ w45781;
	assign w17264 = w17268 ^ w44093;
	assign w17267 = w44097 ^ w17264;
	assign w17364 = w17266 ^ w17267;
	assign w17263 = w17259 ^ w17264;
	assign w17363 = w17262 ^ w17263;
	assign w45366 = ~w17363;
	assign w8599 = w45366 ^ w49704;
	assign w8541 = w8804 ^ w45366;
	assign w8884 = w8541 ^ w8542;
	assign w8819 = w45374 ^ w45366;
	assign w45367 = ~w17364;
	assign w8556 = w45367 ^ w45775;
	assign w8839 = w45375 ^ w45367;
	assign w17493 = w47021 ^ w47027;
	assign w17474 = w17493 & w17478;
	assign w17408 = w17474 ^ w17404;
	assign w17425 = w17426 ^ w17408;
	assign w17382 = w17408 ^ w44099;
	assign w17466 = w17382 ^ w17407;
	assign w17467 = w17473 ^ w17425;
	assign w17464 = w17468 & w17467;
	assign w17459 = w17464 ^ w17424;
	assign w17458 = w17459 & w17460;
	assign w17376 = w17458 ^ w17475;
	assign w17457 = w17458 ^ w17466;
	assign w17434 = w17457 & w17489;
	assign w17443 = w17457 & w47028;
	assign w17463 = w17464 ^ w17466;
	assign w17462 = w17465 & w17463;
	assign w17461 = w17462 ^ w17424;
	assign w17440 = w17461 & w17480;
	assign w17431 = w17461 & w17487;
	assign w17373 = w17462 ^ w17474;
	assign w17370 = w17462 ^ w17418;
	assign w17456 = w17464 ^ w17458;
	assign w17455 = w17466 & w17456;
	assign w17453 = w17455 ^ w17463;
	assign w17452 = w17461 & w17453;
	assign w17375 = w17452 ^ w17476;
	assign w17417 = w17452 ^ w17427;
	assign w17448 = w17417 ^ w17370;
	assign w17433 = w17448 & w17493;
	assign w17451 = w17417 ^ w17419;
	assign w17441 = w17451 & w17490;
	assign w17432 = w17451 & w17486;
	assign w17384 = w17440 ^ w17441;
	assign w17402 = w17440 ^ w17432;
	assign w17442 = w17448 & w17478;
	assign w17400 = w17442 ^ w17433;
	assign w44100 = w17441 ^ w17442;
	assign w44102 = w17455 ^ w17473;
	assign w17414 = w47027 ^ w44102;
	assign w17367 = w17414 ^ w17375;
	assign w17374 = w17404 ^ w17367;
	assign w17447 = w44102 ^ w17425;
	assign w17436 = w17447 & w17488;
	assign w17445 = w17447 & w17484;
	assign w44101 = w17443 ^ w17445;
	assign w17371 = w17376 ^ w17472;
	assign w17450 = w17371 ^ w17374;
	assign w17437 = w17450 & w17482;
	assign w17428 = w17450 & w17491;
	assign w17415 = w17433 ^ w17437;
	assign w17393 = ~w17415;
	assign w17369 = w17373 ^ w17409;
	assign w17372 = w47021 ^ w17369;
	assign w17368 = w47023 ^ w17369;
	assign w17449 = w17371 ^ w17372;
	assign w17439 = w17449 & w17481;
	assign w17430 = w17449 & w17492;
	assign w17394 = w17439 ^ w17428;
	assign w17390 = ~w17394;
	assign w17446 = w17367 ^ w17368;
	assign w17438 = w17446 & w17479;
	assign w17399 = w17438 ^ w17441;
	assign w17429 = w17446 & w17494;
	assign w17396 = ~w17399;
	assign w17423 = w17438 ^ w44100;
	assign w17383 = w17439 ^ w17423;
	assign w17395 = w17438 ^ w17439;
	assign w17389 = w17434 ^ w17423;
	assign w17386 = ~w17389;
	assign w43547 = w17429 ^ w17430;
	assign w17398 = w17402 ^ w43547;
	assign w17397 = w17393 ^ w17398;
	assign w17497 = w17396 ^ w17397;
	assign w17401 = w44101 ^ w17398;
	assign w17498 = w17400 ^ w17401;
	assign w17377 = w17458 ^ w17422;
	assign w17454 = w17414 ^ w17377;
	assign w17435 = w17454 & w17485;
	assign w17444 = w17454 & w17483;
	assign w17411 = w17435 ^ w43547;
	assign w17412 = w17436 ^ w17411;
	assign w49683 = w17412 ^ w17383;
	assign w8799 = w49683 ^ w49698;
	assign w8572 = w8799 ^ w49696;
	assign w8568 = ~w8799;
	assign w8569 = w8568 ^ w49695;
	assign w8566 = w8568 ^ w45526;
	assign w8655 = w8853 ^ w8799;
	assign w17416 = w17444 ^ w17412;
	assign w17385 = w17443 ^ w17416;
	assign w49681 = w17384 ^ w17385;
	assign w17421 = w17445 ^ w17416;
	assign w49682 = w44100 ^ w17421;
	assign w17496 = w17421 ^ w17395;
	assign w45370 = ~w17497;
	assign w45371 = ~w17498;
	assign w45377 = ~w17496;
	assign w17392 = w17393 ^ w17431;
	assign w17388 = w17392 ^ w44101;
	assign w17391 = w17430 ^ w17388;
	assign w17495 = w17390 ^ w17391;
	assign w17387 = w17411 ^ w17388;
	assign w49680 = w17386 ^ w17387;
	assign w45376 = ~w17495;
	assign w45931 = ~w8452;
	assign w8397 = w45931 ^ w49444;
	assign w49326 = w8396 ^ w8397;
	assign w47112 = w49326 ^ w1831;
	assign w12536 = w47114 ^ w47112;
	assign w12521 = w12446 ^ w12536;
	assign w12512 = w12536 & w12521;
	assign w12448 = w47112 ^ w47110;
	assign w12407 = w12448 ^ w47111;
	assign w12531 = w47116 ^ w12407;
	assign w12517 = w47116 & w12531;
	assign w12534 = w47112 ^ w47109;
	assign w12408 = w12448 ^ w12446;
	assign w8240 = w45931 ^ w45780;
	assign w8522 = w8240 ^ w8241;
	assign w49323 = w8522 ^ w8514;
	assign w47115 = w49323 ^ w1828;
	assign w12535 = w47109 ^ w47115;
	assign w12462 = w47115 ^ w47114;
	assign w12445 = w47115 ^ w47113;
	assign w12524 = w12445 ^ w12408;
	assign w12511 = w12533 & w12524;
	assign w12526 = w12445 ^ w12534;
	assign w12525 = w47116 ^ w12526;
	assign w12447 = w47114 ^ w12445;
	assign w12522 = w12452 ^ w12447;
	assign w12523 = w47110 ^ w12447;
	assign w12513 = w12534 & w12523;
	assign w12520 = w47111 ^ w12447;
	assign w12516 = w12535 & w12520;
	assign w12527 = w12462 ^ w12529;
	assign w12518 = w12527 & w12525;
	assign w12449 = w12513 ^ w12447;
	assign w12450 = w12516 ^ w12446;
	assign w12528 = w47115 ^ w12532;
	assign w12515 = w12532 & w12528;
	assign w12530 = w12534 ^ w12462;
	assign w12519 = w12526 & w12530;
	assign w12451 = w12519 ^ w12448;
	assign w12455 = w12451 ^ w12449;
	assign w12460 = w47109 ^ w12455;
	assign w12469 = w12512 ^ w12518;
	assign w12510 = w12469 ^ w12460;
	assign w43891 = w12511 ^ w12517;
	assign w12423 = w12455 ^ w43891;
	assign w12466 = w47111 ^ w12423;
	assign w12461 = w43891 ^ w12446;
	assign w12507 = w12469 ^ w12461;
	assign w8376 = w45931 ^ w49461;
	assign w49337 = w8376 ^ w8377;
	assign w47101 = w49337 ^ w1842;
	assign w27588 = w47103 ^ w47101;
	assign w27663 = w27588 ^ w27678;
	assign w27676 = w47104 ^ w47101;
	assign w27672 = w27676 ^ w27604;
	assign w27671 = w27588 ^ w27594;
	assign w27669 = w27604 ^ w27671;
	assign w27668 = w27587 ^ w27676;
	assign w27667 = w47108 ^ w27668;
	assign w27550 = w27590 ^ w27588;
	assign w27666 = w27587 ^ w27550;
	assign w27677 = w47101 ^ w47107;
	assign w27675 = w47101 ^ w47106;
	assign w27661 = w27668 & w27672;
	assign w27593 = w27661 ^ w27590;
	assign w27660 = w27669 & w27667;
	assign w27658 = w27677 & w27662;
	assign w27592 = w27658 ^ w27588;
	assign w27656 = w27671 & w27664;
	assign w27655 = w27676 & w27665;
	assign w27591 = w27655 ^ w27589;
	assign w27597 = w27593 ^ w27591;
	assign w27602 = w47101 ^ w27597;
	assign w27654 = w27678 & w27663;
	assign w27611 = w27654 ^ w27660;
	assign w27652 = w27611 ^ w27602;
	assign w27563 = w27654 ^ w27655;
	assign w27610 = w27563 ^ w27564;
	assign w27609 = w27610 ^ w27592;
	assign w27651 = w27657 ^ w27609;
	assign w27653 = w27675 & w27666;
	assign w27648 = w27652 & w27651;
	assign w44523 = w27653 ^ w27659;
	assign w27603 = w44523 ^ w27588;
	assign w27649 = w27611 ^ w27603;
	assign w27565 = w27597 ^ w44523;
	assign w27608 = w47103 ^ w27565;
	assign w27643 = w27648 ^ w27608;
	assign w44524 = w27653 ^ w27656;
	assign w27606 = w27654 ^ w44524;
	assign w27562 = w27657 ^ w27606;
	assign w27644 = w47107 ^ w27562;
	assign w27642 = w27643 & w27644;
	assign w27561 = w27642 ^ w27606;
	assign w27560 = w27642 ^ w27659;
	assign w27555 = w27560 ^ w27656;
	assign w27640 = w27648 ^ w27642;
	assign w27566 = w27592 ^ w44524;
	assign w27650 = w27566 ^ w27591;
	assign w27641 = w27642 ^ w27650;
	assign w27647 = w27648 ^ w27650;
	assign w27646 = w27649 & w27647;
	assign w27645 = w27646 ^ w27608;
	assign w27557 = w27646 ^ w27658;
	assign w27553 = w27557 ^ w27593;
	assign w27556 = w47101 ^ w27553;
	assign w27633 = w27555 ^ w27556;
	assign w27554 = w27646 ^ w27602;
	assign w27552 = w47103 ^ w27553;
	assign w27639 = w27650 & w27640;
	assign w27637 = w27639 ^ w27647;
	assign w27636 = w27645 & w27637;
	assign w27601 = w27636 ^ w27611;
	assign w27635 = w27601 ^ w27603;
	assign w27559 = w27636 ^ w27660;
	assign w27632 = w27601 ^ w27554;
	assign w27627 = w27641 & w47108;
	assign w27626 = w27632 & w27662;
	assign w27625 = w27635 & w27674;
	assign w27624 = w27645 & w27664;
	assign w27568 = w27624 ^ w27625;
	assign w27623 = w27633 & w27665;
	assign w27618 = w27641 & w27673;
	assign w27617 = w27632 & w27677;
	assign w27584 = w27626 ^ w27617;
	assign w27616 = w27635 & w27670;
	assign w27586 = w27624 ^ w27616;
	assign w27615 = w27645 & w27671;
	assign w27614 = w27633 & w27676;
	assign w44525 = w27625 ^ w27626;
	assign w44527 = w27639 ^ w27657;
	assign w27598 = w47107 ^ w44527;
	assign w27638 = w27598 ^ w27561;
	assign w27619 = w27638 & w27669;
	assign w27628 = w27638 & w27667;
	assign w27551 = w27598 ^ w27559;
	assign w27558 = w27588 ^ w27551;
	assign w27634 = w27555 ^ w27558;
	assign w27621 = w27634 & w27666;
	assign w27599 = w27617 ^ w27621;
	assign w27577 = ~w27599;
	assign w27576 = w27577 ^ w27615;
	assign w27630 = w27551 ^ w27552;
	assign w27613 = w27630 & w27678;
	assign w27612 = w27634 & w27675;
	assign w27578 = w27623 ^ w27612;
	assign w27574 = ~w27578;
	assign w43578 = w27613 ^ w27614;
	assign w27595 = w27619 ^ w43578;
	assign w27582 = w27586 ^ w43578;
	assign w27581 = w27577 ^ w27582;
	assign w27622 = w27630 & w27663;
	assign w27579 = w27622 ^ w27623;
	assign w27607 = w27622 ^ w44525;
	assign w27573 = w27618 ^ w27607;
	assign w27570 = ~w27573;
	assign w27567 = w27623 ^ w27607;
	assign w27583 = w27622 ^ w27625;
	assign w27580 = ~w27583;
	assign w27681 = w27580 ^ w27581;
	assign w27631 = w44527 ^ w27609;
	assign w27629 = w27631 & w27668;
	assign w27620 = w27631 & w27672;
	assign w27596 = w27620 ^ w27595;
	assign w27600 = w27628 ^ w27596;
	assign w27605 = w27629 ^ w27600;
	assign w49674 = w44525 ^ w27605;
	assign w27680 = w27605 ^ w27579;
	assign w27569 = w27627 ^ w27600;
	assign w49673 = w27568 ^ w27569;
	assign w49675 = w27596 ^ w27567;
	assign w8813 = w49674 ^ w49678;
	assign w8800 = w49671 ^ w49675;
	assign w8792 = w49675 ^ w49679;
	assign w8701 = w8811 ^ w8792;
	assign w49554 = w49671 ^ w8701;
	assign w49551 = w8879 ^ w8813;
	assign w8559 = w8800 ^ w45705;
	assign w8564 = w49673 ^ w8552;
	assign w8565 = ~w8800;
	assign w8563 = w8565 ^ w49678;
	assign w8874 = w8563 ^ w8564;
	assign w49567 = w8874 ^ w8821;
	assign w46944 = w49567 ^ w915;
	assign w8662 = ~w49674;
	assign w8683 = w8792 ^ w45242;
	assign w8659 = w8817 ^ w8813;
	assign w8687 = w8689 ^ w8813;
	assign w8668 = w8792 ^ w49673;
	assign w8672 = w8833 ^ w8792;
	assign w8677 = w8662 ^ w49670;
	assign w49568 = w8676 ^ w8677;
	assign w8661 = w8792 ^ w8662;
	assign w49562 = w8683 ^ w8684;
	assign w46960 = w49551 ^ w899;
	assign w46957 = w49554 ^ w902;
	assign w27408 = w46960 ^ w46957;
	assign w46949 = w49562 ^ w910;
	assign w46943 = w49568 ^ w916;
	assign w8818 = w49673 ^ w49677;
	assign w8690 = w8681 ^ w8818;
	assign w49550 = w8880 ^ w8818;
	assign w8660 = w8663 ^ w8818;
	assign w49575 = w8660 ^ w8661;
	assign w46936 = w49575 ^ w923;
	assign w46961 = w49550 ^ w898;
	assign w44526 = w27627 ^ w27629;
	assign w27585 = w44526 ^ w27582;
	assign w27682 = w27584 ^ w27585;
	assign w27572 = w27576 ^ w44526;
	assign w27575 = w27614 ^ w27572;
	assign w27679 = w27574 ^ w27575;
	assign w27571 = w27595 ^ w27572;
	assign w49672 = w27570 ^ w27571;
	assign w8823 = w49672 ^ w49676;
	assign w8562 = w49672 ^ w49668;
	assign w8692 = w8832 ^ w8823;
	assign w49557 = w49663 ^ w8692;
	assign w8667 = w8825 ^ w8823;
	assign w49574 = w8667 ^ w8668;
	assign w8706 = w8823 ^ w45705;
	assign w49549 = w8706 ^ w8707;
	assign w46962 = w49549 ^ w897;
	assign w27410 = w46962 ^ w46960;
	assign w27296 = w46961 ^ w46962;
	assign w27407 = w46957 ^ w46962;
	assign w46937 = w49574 ^ w922;
	assign w46954 = w49557 ^ w905;
	assign w8561 = w8800 ^ w49677;
	assign w8875 = w8561 ^ w8562;
	assign w49566 = w8875 ^ w8825;
	assign w46945 = w49566 ^ w914;
	assign w8682 = w8833 ^ w8800;
	assign w49563 = w45698 ^ w8682;
	assign w46948 = w49563 ^ w911;
	assign w12131 = w46949 ^ w46954;
	assign w45618 = ~w27680;
	assign w8810 = w45242 ^ w45618;
	assign w8657 = w49675 ^ w45618;
	assign w49578 = w8656 ^ w8657;
	assign w46933 = w49578 ^ w926;
	assign w8673 = w8810 ^ w8793;
	assign w49570 = w49679 ^ w8673;
	assign w49561 = w45618 ^ w8685;
	assign w46950 = w49561 ^ w909;
	assign w8702 = w8810 ^ w45704;
	assign w46941 = w49570 ^ w918;
	assign w16956 = w46944 ^ w46941;
	assign w16868 = w46943 ^ w46941;
	assign w24192 = w46936 ^ w46933;
	assign w49553 = w8702 ^ w8703;
	assign w46958 = w49553 ^ w901;
	assign w27322 = w46960 ^ w46958;
	assign w45619 = ~w27681;
	assign w8826 = w45619 ^ w45705;
	assign w49548 = w8881 ^ w8826;
	assign w8671 = w8792 ^ w45619;
	assign w8669 = w8828 ^ w8826;
	assign w49573 = w49672 ^ w8669;
	assign w8680 = w45619 ^ w12271;
	assign w49565 = w8679 ^ w8680;
	assign w8694 = w8833 ^ w8826;
	assign w46963 = w49548 ^ w896;
	assign w27319 = w46963 ^ w46961;
	assign w27321 = w46962 ^ w27319;
	assign w27397 = w46958 ^ w27321;
	assign w27400 = w27319 ^ w27408;
	assign w27336 = w46963 ^ w46962;
	assign w27404 = w27408 ^ w27336;
	assign w27409 = w46957 ^ w46963;
	assign w27393 = w27400 & w27404;
	assign w27325 = w27393 ^ w27322;
	assign w27387 = w27408 & w27397;
	assign w27323 = w27387 ^ w27321;
	assign w27329 = w27325 ^ w27323;
	assign w27334 = w46957 ^ w27329;
	assign w46938 = w49573 ^ w921;
	assign w24191 = w46933 ^ w46938;
	assign w46946 = w49565 ^ w913;
	assign w16844 = w46945 ^ w46946;
	assign w16958 = w46946 ^ w46944;
	assign w16943 = w16868 ^ w16958;
	assign w16934 = w16958 & w16943;
	assign w24080 = w46937 ^ w46938;
	assign w24194 = w46938 ^ w46936;
	assign w16955 = w46941 ^ w46946;
	assign w45620 = ~w27682;
	assign w8830 = w45620 ^ w45698;
	assign w8696 = w8830 ^ w8793;
	assign w49555 = w45616 ^ w8696;
	assign w8560 = w45620 ^ w45243;
	assign w8876 = w8559 ^ w8560;
	assign w8670 = w8832 ^ w8830;
	assign w49572 = w8670 ^ w8671;
	assign w49571 = w45620 ^ w8672;
	assign w46939 = w49572 ^ w920;
	assign w24193 = w46933 ^ w46939;
	assign w24120 = w46939 ^ w46938;
	assign w46940 = w49571 ^ w919;
	assign w8708 = w8830 ^ w8802;
	assign w49547 = w45243 ^ w8708;
	assign w46964 = w49547 ^ w895;
	assign w27399 = w46964 ^ w27400;
	assign w27326 = w46964 ^ w46958;
	assign w27396 = w27326 ^ w27321;
	assign w46956 = w49555 ^ w903;
	assign w12050 = w46956 ^ w46950;
	assign w24188 = w24192 ^ w24120;
	assign w24103 = w46939 ^ w46937;
	assign w24105 = w46938 ^ w24103;
	assign w24184 = w24103 ^ w24192;
	assign w24177 = w24184 & w24188;
	assign w24183 = w46940 ^ w24184;
	assign w49564 = w8876 ^ w8832;
	assign w46947 = w49564 ^ w912;
	assign w16867 = w46947 ^ w46945;
	assign w16948 = w16867 ^ w16956;
	assign w16884 = w46947 ^ w46946;
	assign w16869 = w46946 ^ w16867;
	assign w16947 = w46948 ^ w16948;
	assign w16952 = w16956 ^ w16884;
	assign w16941 = w16948 & w16952;
	assign w16957 = w46941 ^ w46947;
	assign w16942 = w46943 ^ w16869;
	assign w16938 = w16957 & w16942;
	assign w16872 = w16938 ^ w16868;
	assign w45625 = ~w27679;
	assign w49576 = w45625 ^ w8659;
	assign w8674 = w8811 ^ w45625;
	assign w49569 = w8674 ^ w8675;
	assign w46942 = w49569 ^ w917;
	assign w16870 = w46944 ^ w46942;
	assign w16873 = w16941 ^ w16870;
	assign w16874 = w46948 ^ w46942;
	assign w16951 = w16868 ^ w16874;
	assign w16954 = w46943 ^ w16874;
	assign w16949 = w16884 ^ w16951;
	assign w16940 = w16949 & w16947;
	assign w16944 = w16874 ^ w16869;
	assign w16891 = w16934 ^ w16940;
	assign w16950 = w46947 ^ w16954;
	assign w16937 = w16954 & w16950;
	assign w16945 = w46942 ^ w16869;
	assign w46935 = w49576 ^ w924;
	assign w24178 = w46935 ^ w24105;
	assign w24174 = w24193 & w24178;
	assign w16936 = w16951 & w16944;
	assign w16935 = w16956 & w16945;
	assign w16843 = w16934 ^ w16935;
	assign w16890 = w16843 ^ w16844;
	assign w16889 = w16890 ^ w16872;
	assign w16931 = w16937 ^ w16889;
	assign w16871 = w16935 ^ w16869;
	assign w16877 = w16873 ^ w16871;
	assign w16882 = w46941 ^ w16877;
	assign w16932 = w16891 ^ w16882;
	assign w16830 = w16870 ^ w16868;
	assign w16928 = w16932 & w16931;
	assign w16946 = w16867 ^ w16830;
	assign w16933 = w16955 & w16946;
	assign w8808 = w45625 ^ w45703;
	assign w8686 = w8821 ^ w8808;
	assign w49560 = w45621 ^ w8686;
	assign w8658 = w8810 ^ w8808;
	assign w49577 = w45614 ^ w8658;
	assign w46934 = w49577 ^ w925;
	assign w24110 = w46940 ^ w46934;
	assign w24106 = w46936 ^ w46934;
	assign w24065 = w24106 ^ w46935;
	assign w24189 = w46940 ^ w24065;
	assign w24109 = w24177 ^ w24106;
	assign w24175 = w46940 & w24189;
	assign w24190 = w46935 ^ w24110;
	assign w24186 = w46939 ^ w24190;
	assign w24173 = w24190 & w24186;
	assign w24181 = w46934 ^ w24105;
	assign w24171 = w24192 & w24181;
	assign w24107 = w24171 ^ w24105;
	assign w24113 = w24109 ^ w24107;
	assign w24118 = w46933 ^ w24113;
	assign w46951 = w49560 ^ w908;
	assign w12130 = w46951 ^ w12050;
	assign w12044 = w46951 ^ w46949;
	assign w12127 = w12044 ^ w12050;
	assign w8704 = w8808 ^ w49678;
	assign w24180 = w24110 ^ w24105;
	assign w49552 = w8704 ^ w8705;
	assign w46959 = w49552 ^ w900;
	assign w27394 = w46959 ^ w27321;
	assign w27320 = w46959 ^ w46957;
	assign w27395 = w27320 ^ w27410;
	assign w27403 = w27320 ^ w27326;
	assign w27401 = w27336 ^ w27403;
	assign w27406 = w46959 ^ w27326;
	assign w27402 = w46963 ^ w27406;
	assign w27282 = w27322 ^ w27320;
	assign w27398 = w27319 ^ w27282;
	assign w27281 = w27322 ^ w46959;
	assign w27405 = w46964 ^ w27281;
	assign w27392 = w27401 & w27399;
	assign w27391 = w46964 & w27405;
	assign w27390 = w27409 & w27394;
	assign w27324 = w27390 ^ w27320;
	assign w27389 = w27406 & w27402;
	assign w27388 = w27403 & w27396;
	assign w27386 = w27410 & w27395;
	assign w27343 = w27386 ^ w27392;
	assign w27384 = w27343 ^ w27334;
	assign w27295 = w27386 ^ w27387;
	assign w27342 = w27295 ^ w27296;
	assign w27341 = w27342 ^ w27324;
	assign w27383 = w27389 ^ w27341;
	assign w27385 = w27407 & w27398;
	assign w27380 = w27384 & w27383;
	assign w44077 = w16933 ^ w16936;
	assign w16886 = w16934 ^ w44077;
	assign w16842 = w16937 ^ w16886;
	assign w16924 = w46947 ^ w16842;
	assign w16846 = w16872 ^ w44077;
	assign w16930 = w16846 ^ w16871;
	assign w16927 = w16928 ^ w16930;
	assign w24104 = w46935 ^ w46933;
	assign w24108 = w24174 ^ w24104;
	assign w24066 = w24106 ^ w24104;
	assign w24187 = w24104 ^ w24110;
	assign w24172 = w24187 & w24180;
	assign w24182 = w24103 ^ w24066;
	assign w24169 = w24191 & w24182;
	assign w24185 = w24120 ^ w24187;
	assign w24176 = w24185 & w24183;
	assign w24179 = w24104 ^ w24194;
	assign w24170 = w24194 & w24179;
	assign w24079 = w24170 ^ w24171;
	assign w24126 = w24079 ^ w24080;
	assign w24125 = w24126 ^ w24108;
	assign w24127 = w24170 ^ w24176;
	assign w24167 = w24173 ^ w24125;
	assign w44380 = w24169 ^ w24175;
	assign w24119 = w44380 ^ w24104;
	assign w24165 = w24127 ^ w24119;
	assign w24081 = w24113 ^ w44380;
	assign w24124 = w46935 ^ w24081;
	assign w44381 = w24169 ^ w24172;
	assign w24122 = w24170 ^ w44381;
	assign w24078 = w24173 ^ w24122;
	assign w24160 = w46939 ^ w24078;
	assign w24082 = w24108 ^ w44381;
	assign w24166 = w24082 ^ w24107;
	assign w24168 = w24127 ^ w24118;
	assign w24164 = w24168 & w24167;
	assign w24163 = w24164 ^ w24166;
	assign w24162 = w24165 & w24163;
	assign w24073 = w24162 ^ w24174;
	assign w24069 = w24073 ^ w24109;
	assign w24070 = w24162 ^ w24118;
	assign w24072 = w46933 ^ w24069;
	assign w24068 = w46935 ^ w24069;
	assign w24159 = w24164 ^ w24124;
	assign w24158 = w24159 & w24160;
	assign w24077 = w24158 ^ w24122;
	assign w24156 = w24164 ^ w24158;
	assign w24155 = w24166 & w24156;
	assign w24157 = w24158 ^ w24166;
	assign w24143 = w24157 & w46940;
	assign w24076 = w24158 ^ w24175;
	assign w24134 = w24157 & w24189;
	assign w24153 = w24155 ^ w24163;
	assign w24071 = w24076 ^ w24172;
	assign w24149 = w24071 ^ w24072;
	assign w24139 = w24149 & w24181;
	assign w24130 = w24149 & w24192;
	assign w44384 = w24155 ^ w24173;
	assign w24114 = w46939 ^ w44384;
	assign w24154 = w24114 ^ w24077;
	assign w24144 = w24154 & w24183;
	assign w24135 = w24154 & w24185;
	assign w24147 = w44384 ^ w24125;
	assign w24145 = w24147 & w24184;
	assign w24136 = w24147 & w24188;
	assign w44383 = w24143 ^ w24145;
	assign w44512 = w27385 ^ w27388;
	assign w27298 = w27324 ^ w44512;
	assign w27382 = w27298 ^ w27323;
	assign w27379 = w27380 ^ w27382;
	assign w27338 = w27386 ^ w44512;
	assign w27294 = w27389 ^ w27338;
	assign w27376 = w46963 ^ w27294;
	assign w44515 = w27385 ^ w27391;
	assign w27297 = w27329 ^ w44515;
	assign w27340 = w46959 ^ w27297;
	assign w27375 = w27380 ^ w27340;
	assign w27374 = w27375 & w27376;
	assign w27372 = w27380 ^ w27374;
	assign w27293 = w27374 ^ w27338;
	assign w27292 = w27374 ^ w27391;
	assign w27287 = w27292 ^ w27388;
	assign w27371 = w27382 & w27372;
	assign w27369 = w27371 ^ w27379;
	assign w44514 = w27371 ^ w27389;
	assign w27363 = w44514 ^ w27341;
	assign w27352 = w27363 & w27404;
	assign w27361 = w27363 & w27400;
	assign w27330 = w46963 ^ w44514;
	assign w27370 = w27330 ^ w27293;
	assign w27360 = w27370 & w27399;
	assign w27351 = w27370 & w27401;
	assign w27373 = w27374 ^ w27382;
	assign w27359 = w27373 & w46964;
	assign w27350 = w27373 & w27405;
	assign w27335 = w44515 ^ w27320;
	assign w27381 = w27343 ^ w27335;
	assign w27378 = w27381 & w27379;
	assign w27377 = w27378 ^ w27340;
	assign w27289 = w27378 ^ w27390;
	assign w27285 = w27289 ^ w27325;
	assign w27288 = w46957 ^ w27285;
	assign w27365 = w27287 ^ w27288;
	assign w27286 = w27378 ^ w27334;
	assign w27284 = w46959 ^ w27285;
	assign w27368 = w27377 & w27369;
	assign w27333 = w27368 ^ w27343;
	assign w27367 = w27333 ^ w27335;
	assign w27291 = w27368 ^ w27392;
	assign w27283 = w27330 ^ w27291;
	assign w27290 = w27320 ^ w27283;
	assign w27366 = w27287 ^ w27290;
	assign w27364 = w27333 ^ w27286;
	assign w27362 = w27283 ^ w27284;
	assign w27358 = w27364 & w27394;
	assign w27357 = w27367 & w27406;
	assign w27356 = w27377 & w27396;
	assign w27300 = w27356 ^ w27357;
	assign w27355 = w27365 & w27397;
	assign w27354 = w27362 & w27395;
	assign w27315 = w27354 ^ w27357;
	assign w27312 = ~w27315;
	assign w27311 = w27354 ^ w27355;
	assign w27353 = w27366 & w27398;
	assign w27349 = w27364 & w27409;
	assign w27331 = w27349 ^ w27353;
	assign w27316 = w27358 ^ w27349;
	assign w27309 = ~w27331;
	assign w27348 = w27367 & w27402;
	assign w27318 = w27356 ^ w27348;
	assign w27347 = w27377 & w27403;
	assign w27308 = w27309 ^ w27347;
	assign w27346 = w27365 & w27408;
	assign w27345 = w27362 & w27410;
	assign w27344 = w27366 & w27407;
	assign w27310 = w27355 ^ w27344;
	assign w27306 = ~w27310;
	assign w44513 = w27345 ^ w27346;
	assign w27327 = w27351 ^ w44513;
	assign w27328 = w27352 ^ w27327;
	assign w27332 = w27360 ^ w27328;
	assign w27301 = w27359 ^ w27332;
	assign w49845 = w27300 ^ w27301;
	assign w27337 = w27361 ^ w27332;
	assign w27412 = w27337 ^ w27311;
	assign w27314 = w27318 ^ w44513;
	assign w27313 = w27309 ^ w27314;
	assign w27413 = w27312 ^ w27313;
	assign w44516 = w27357 ^ w27358;
	assign w49846 = w44516 ^ w27337;
	assign w27339 = w27354 ^ w44516;
	assign w27305 = w27350 ^ w27339;
	assign w27302 = ~w27305;
	assign w27299 = w27355 ^ w27339;
	assign w49847 = w27328 ^ w27299;
	assign w44517 = w27359 ^ w27361;
	assign w27317 = w44517 ^ w27314;
	assign w27414 = w27316 ^ w27317;
	assign w27304 = w27308 ^ w44517;
	assign w27307 = w27346 ^ w27304;
	assign w27411 = w27306 ^ w27307;
	assign w27303 = w27327 ^ w27304;
	assign w49844 = w27302 ^ w27303;
	assign w16829 = w16870 ^ w46943;
	assign w16953 = w46948 ^ w16829;
	assign w16939 = w46948 & w16953;
	assign w44076 = w16933 ^ w16939;
	assign w16883 = w44076 ^ w16868;
	assign w16929 = w16891 ^ w16883;
	assign w16926 = w16929 & w16927;
	assign w16834 = w16926 ^ w16882;
	assign w16837 = w16926 ^ w16938;
	assign w16833 = w16837 ^ w16873;
	assign w16832 = w46943 ^ w16833;
	assign w16836 = w46941 ^ w16833;
	assign w16845 = w16877 ^ w44076;
	assign w16888 = w46943 ^ w16845;
	assign w16923 = w16928 ^ w16888;
	assign w16925 = w16926 ^ w16888;
	assign w16922 = w16923 & w16924;
	assign w16921 = w16922 ^ w16930;
	assign w16907 = w16921 & w46948;
	assign w16840 = w16922 ^ w16939;
	assign w16835 = w16840 ^ w16936;
	assign w16920 = w16928 ^ w16922;
	assign w16898 = w16921 & w16953;
	assign w16913 = w16835 ^ w16836;
	assign w16894 = w16913 & w16956;
	assign w16903 = w16913 & w16945;
	assign w16919 = w16930 & w16920;
	assign w16917 = w16919 ^ w16927;
	assign w16916 = w16925 & w16917;
	assign w16839 = w16916 ^ w16940;
	assign w16881 = w16916 ^ w16891;
	assign w16915 = w16881 ^ w16883;
	assign w16896 = w16915 & w16950;
	assign w16912 = w16881 ^ w16834;
	assign w16905 = w16915 & w16954;
	assign w44080 = w16919 ^ w16937;
	assign w16878 = w46947 ^ w44080;
	assign w16831 = w16878 ^ w16839;
	assign w16910 = w16831 ^ w16832;
	assign w16838 = w16868 ^ w16831;
	assign w16914 = w16835 ^ w16838;
	assign w16901 = w16914 & w16946;
	assign w16892 = w16914 & w16955;
	assign w16858 = w16903 ^ w16892;
	assign w16854 = ~w16858;
	assign w16911 = w44080 ^ w16889;
	assign w16900 = w16911 & w16952;
	assign w16909 = w16911 & w16948;
	assign w44079 = w16907 ^ w16909;
	assign w16906 = w16912 & w16942;
	assign w44078 = w16905 ^ w16906;
	assign w16841 = w16922 ^ w16886;
	assign w16918 = w16878 ^ w16841;
	assign w16908 = w16918 & w16947;
	assign w16904 = w16925 & w16944;
	assign w16866 = w16904 ^ w16896;
	assign w16848 = w16904 ^ w16905;
	assign w16902 = w16910 & w16943;
	assign w16887 = w16902 ^ w44078;
	assign w16853 = w16898 ^ w16887;
	assign w16859 = w16902 ^ w16903;
	assign w16863 = w16902 ^ w16905;
	assign w16850 = ~w16853;
	assign w16847 = w16903 ^ w16887;
	assign w16860 = ~w16863;
	assign w16899 = w16918 & w16949;
	assign w16897 = w16912 & w16957;
	assign w16879 = w16897 ^ w16901;
	assign w16864 = w16906 ^ w16897;
	assign w16857 = ~w16879;
	assign w16895 = w16925 & w16951;
	assign w16856 = w16857 ^ w16895;
	assign w16852 = w16856 ^ w44079;
	assign w16855 = w16894 ^ w16852;
	assign w16959 = w16854 ^ w16855;
	assign w45359 = ~w16959;
	assign w16893 = w16910 & w16958;
	assign w43545 = w16893 ^ w16894;
	assign w16875 = w16899 ^ w43545;
	assign w16851 = w16875 ^ w16852;
	assign w49892 = w16850 ^ w16851;
	assign w16876 = w16900 ^ w16875;
	assign w16880 = w16908 ^ w16876;
	assign w16849 = w16907 ^ w16880;
	assign w16885 = w16909 ^ w16880;
	assign w16960 = w16885 ^ w16859;
	assign w49893 = w16848 ^ w16849;
	assign w49895 = w16876 ^ w16847;
	assign w49894 = w44078 ^ w16885;
	assign w16862 = w16866 ^ w43545;
	assign w16861 = w16857 ^ w16862;
	assign w16865 = w44079 ^ w16862;
	assign w16962 = w16864 ^ w16865;
	assign w16961 = w16860 ^ w16861;
	assign w45354 = ~w16962;
	assign w45360 = ~w16960;
	assign w45361 = ~w16961;
	assign w45610 = ~w27412;
	assign w45611 = ~w27413;
	assign w45612 = ~w27414;
	assign w45617 = ~w27411;
	assign w24161 = w24162 ^ w24124;
	assign w24140 = w24161 & w24180;
	assign w24152 = w24161 & w24153;
	assign w24131 = w24161 & w24187;
	assign w24117 = w24152 ^ w24127;
	assign w24148 = w24117 ^ w24070;
	assign w24133 = w24148 & w24193;
	assign w24142 = w24148 & w24178;
	assign w24075 = w24152 ^ w24176;
	assign w24100 = w24142 ^ w24133;
	assign w24151 = w24117 ^ w24119;
	assign w24132 = w24151 & w24186;
	assign w24141 = w24151 & w24190;
	assign w24084 = w24140 ^ w24141;
	assign w24102 = w24140 ^ w24132;
	assign w24067 = w24114 ^ w24075;
	assign w24074 = w24104 ^ w24067;
	assign w24150 = w24071 ^ w24074;
	assign w24137 = w24150 & w24182;
	assign w24146 = w24067 ^ w24068;
	assign w24129 = w24146 & w24194;
	assign w24128 = w24150 & w24191;
	assign w24094 = w24139 ^ w24128;
	assign w43565 = w24129 ^ w24130;
	assign w24098 = w24102 ^ w43565;
	assign w24101 = w44383 ^ w24098;
	assign w24111 = w24135 ^ w43565;
	assign w24112 = w24136 ^ w24111;
	assign w24116 = w24144 ^ w24112;
	assign w24085 = w24143 ^ w24116;
	assign w49878 = w24084 ^ w24085;
	assign w24121 = w24145 ^ w24116;
	assign w24198 = w24100 ^ w24101;
	assign w44382 = w24141 ^ w24142;
	assign w49879 = w44382 ^ w24121;
	assign w24138 = w24146 & w24179;
	assign w24095 = w24138 ^ w24139;
	assign w24196 = w24121 ^ w24095;
	assign w24123 = w24138 ^ w44382;
	assign w24089 = w24134 ^ w24123;
	assign w24083 = w24139 ^ w24123;
	assign w49880 = w24112 ^ w24083;
	assign w24086 = ~w24089;
	assign w24099 = w24138 ^ w24141;
	assign w24096 = ~w24099;
	assign w24115 = w24133 ^ w24137;
	assign w24093 = ~w24115;
	assign w24097 = w24093 ^ w24098;
	assign w24197 = w24096 ^ w24097;
	assign w45523 = ~w24196;
	assign w45524 = ~w24197;
	assign w45525 = ~w24198;
	assign w24090 = ~w24094;
	assign w24092 = w24093 ^ w24131;
	assign w24088 = w24092 ^ w44383;
	assign w24091 = w24130 ^ w24088;
	assign w24087 = w24111 ^ w24088;
	assign w49877 = w24086 ^ w24087;
	assign w12421 = w12512 ^ w12513;
	assign w12468 = w12421 ^ w12422;
	assign w12467 = w12468 ^ w12450;
	assign w12509 = w12515 ^ w12467;
	assign w12506 = w12510 & w12509;
	assign w12501 = w12506 ^ w12466;
	assign w12514 = w12529 & w12522;
	assign w43892 = w12511 ^ w12514;
	assign w12464 = w12512 ^ w43892;
	assign w12420 = w12515 ^ w12464;
	assign w12424 = w12450 ^ w43892;
	assign w12508 = w12424 ^ w12449;
	assign w12505 = w12506 ^ w12508;
	assign w12504 = w12507 & w12505;
	assign w12412 = w12504 ^ w12460;
	assign w12503 = w12504 ^ w12466;
	assign w12473 = w12503 & w12529;
	assign w12482 = w12503 & w12522;
	assign w12415 = w12504 ^ w12516;
	assign w12411 = w12415 ^ w12451;
	assign w12414 = w47109 ^ w12411;
	assign w12410 = w47111 ^ w12411;
	assign w12502 = w47115 ^ w12420;
	assign w12500 = w12501 & w12502;
	assign w12419 = w12500 ^ w12464;
	assign w12499 = w12500 ^ w12508;
	assign w12485 = w12499 & w47116;
	assign w12476 = w12499 & w12531;
	assign w12498 = w12506 ^ w12500;
	assign w12418 = w12500 ^ w12517;
	assign w12413 = w12418 ^ w12514;
	assign w12491 = w12413 ^ w12414;
	assign w12472 = w12491 & w12534;
	assign w12481 = w12491 & w12523;
	assign w12497 = w12508 & w12498;
	assign w12495 = w12497 ^ w12505;
	assign w12494 = w12503 & w12495;
	assign w12459 = w12494 ^ w12469;
	assign w12490 = w12459 ^ w12412;
	assign w12484 = w12490 & w12520;
	assign w12475 = w12490 & w12535;
	assign w12417 = w12494 ^ w12518;
	assign w12493 = w12459 ^ w12461;
	assign w12474 = w12493 & w12528;
	assign w12444 = w12482 ^ w12474;
	assign w12483 = w12493 & w12532;
	assign w12426 = w12482 ^ w12483;
	assign w12442 = w12484 ^ w12475;
	assign w43894 = w12483 ^ w12484;
	assign w43896 = w12497 ^ w12515;
	assign w12489 = w43896 ^ w12467;
	assign w12478 = w12489 & w12530;
	assign w12456 = w47115 ^ w43896;
	assign w12409 = w12456 ^ w12417;
	assign w12416 = w12446 ^ w12409;
	assign w12492 = w12413 ^ w12416;
	assign w12479 = w12492 & w12524;
	assign w12457 = w12475 ^ w12479;
	assign w12435 = ~w12457;
	assign w12434 = w12435 ^ w12473;
	assign w12470 = w12492 & w12533;
	assign w12436 = w12481 ^ w12470;
	assign w12432 = ~w12436;
	assign w12488 = w12409 ^ w12410;
	assign w12471 = w12488 & w12536;
	assign w12480 = w12488 & w12521;
	assign w12437 = w12480 ^ w12481;
	assign w12465 = w12480 ^ w43894;
	assign w12425 = w12481 ^ w12465;
	assign w12431 = w12476 ^ w12465;
	assign w12428 = ~w12431;
	assign w12496 = w12456 ^ w12419;
	assign w12477 = w12496 & w12527;
	assign w12486 = w12496 & w12525;
	assign w12441 = w12480 ^ w12483;
	assign w12438 = ~w12441;
	assign w43893 = w12471 ^ w12472;
	assign w12453 = w12477 ^ w43893;
	assign w12454 = w12478 ^ w12453;
	assign w12458 = w12486 ^ w12454;
	assign w12427 = w12485 ^ w12458;
	assign w49686 = w12426 ^ w12427;
	assign w8842 = w49681 ^ w49686;
	assign w8571 = ~w49686;
	assign w8581 = w49692 ^ w8571;
	assign w8570 = w8571 ^ w49680;
	assign w8872 = w8569 ^ w8570;
	assign w49582 = w8872 ^ w8831;
	assign w8609 = ~w8842;
	assign w8632 = w8609 ^ w8822;
	assign w8607 = w8609 ^ w8841;
	assign w46929 = w49582 ^ w866;
	assign w49690 = w12454 ^ w12425;
	assign w8794 = w49683 ^ w49690;
	assign w8601 = w8805 ^ w8794;
	assign w49610 = w49694 ^ w8601;
	assign w8640 = w8853 ^ w8794;
	assign w49587 = w45371 ^ w8640;
	assign w46924 = w49587 ^ w871;
	assign w8642 = w49690 ^ w45377;
	assign w49586 = w8641 ^ w8642;
	assign w46925 = w49586 ^ w870;
	assign w46901 = w49610 ^ w894;
	assign w8798 = w49690 ^ w49694;
	assign w8579 = ~w8798;
	assign w8580 = w8579 ^ w49697;
	assign w8868 = w8580 ^ w8581;
	assign w8574 = w8798 ^ w45533;
	assign w8576 = w8579 ^ w49696;
	assign w12440 = w12444 ^ w43893;
	assign w12487 = w12489 & w12526;
	assign w12463 = w12487 ^ w12458;
	assign w12538 = w12463 ^ w12437;
	assign w49689 = ~w12538;
	assign w8820 = w45377 ^ w49689;
	assign w8617 = w45385 ^ w12538;
	assign w8602 = w8820 ^ w8816;
	assign w49609 = w45385 ^ w8602;
	assign w8645 = w12538 ^ w45376;
	assign w8643 = w8644 ^ w8645;
	assign w8620 = w8820 ^ w45532;
	assign w49585 = ~w8643;
	assign w8618 = ~w8620;
	assign w46902 = w49609 ^ w893;
	assign w49687 = w43894 ^ w12463;
	assign w8834 = w49682 ^ w49687;
	assign w49599 = w8868 ^ w8834;
	assign w8573 = w49687 ^ w49681;
	assign w8871 = w8572 ^ w8573;
	assign w49583 = w8871 ^ w8822;
	assign w8622 = w49693 ^ w49687;
	assign w8631 = w8834 ^ w8816;
	assign w49592 = w45376 ^ w8631;
	assign w46928 = w49583 ^ w867;
	assign w16822 = w46928 ^ w46925;
	assign w46912 = w49599 ^ w883;
	assign w46926 = w49585 ^ w869;
	assign w16736 = w46928 ^ w46926;
	assign w8606 = ~w8834;
	assign w8604 = w8606 ^ w8831;
	assign w8629 = w8820 ^ w8791;
	assign w49594 = w49683 ^ w8629;
	assign w46917 = w49594 ^ w878;
	assign w43895 = w12485 ^ w12487;
	assign w12443 = w43895 ^ w12440;
	assign w12540 = w12442 ^ w12443;
	assign w12430 = w12434 ^ w43895;
	assign w12433 = w12472 ^ w12430;
	assign w12429 = w12453 ^ w12430;
	assign w12537 = w12432 ^ w12433;
	assign w49688 = ~w12537;
	assign w8650 = w12537 ^ w49682;
	assign w49584 = w8649 ^ w8650;
	assign w8619 = w45384 ^ w12537;
	assign w46927 = w49584 ^ w868;
	assign w16734 = w46927 ^ w46925;
	assign w16696 = w16736 ^ w16734;
	assign w49685 = w12428 ^ w12429;
	assign w8849 = w49680 ^ w49685;
	assign w8578 = ~w49685;
	assign w8577 = w49691 ^ w8578;
	assign w8869 = w8576 ^ w8577;
	assign w8653 = w8578 ^ w45370;
	assign w49581 = w8652 ^ w8653;
	assign w8610 = w8849 ^ w8845;
	assign w49605 = w49691 ^ w8610;
	assign w49598 = w8869 ^ w8842;
	assign w46913 = w49598 ^ w882;
	assign w49601 = w8618 ^ w8619;
	assign w46910 = w49601 ^ w885;
	assign w27188 = w46912 ^ w46910;
	assign w46930 = w49581 ^ w865;
	assign w16710 = w46929 ^ w46930;
	assign w16821 = w46925 ^ w46930;
	assign w16824 = w46930 ^ w46928;
	assign w16809 = w16734 ^ w16824;
	assign w16800 = w16824 & w16809;
	assign w8625 = ~w8849;
	assign w8634 = w8625 ^ w8831;
	assign w8623 = w8625 ^ w49695;
	assign w46906 = w49605 ^ w889;
	assign w30355 = w46901 ^ w46906;
	assign w8827 = w45376 ^ w49688;
	assign w8603 = w8827 ^ w8822;
	assign w49608 = w45384 ^ w8603;
	assign w8621 = w8827 ^ w45531;
	assign w49600 = w8621 ^ w8622;
	assign w46911 = w49600 ^ w884;
	assign w27147 = w27188 ^ w46911;
	assign w8630 = w8827 ^ w8805;
	assign w49593 = w45377 ^ w8630;
	assign w46918 = w49593 ^ w877;
	assign w11916 = w46924 ^ w46918;
	assign w46903 = w49608 ^ w892;
	assign w30268 = w46903 ^ w46901;
	assign w46919 = w49592 ^ w876;
	assign w11910 = w46919 ^ w46917;
	assign w11993 = w11910 ^ w11916;
	assign w45246 = ~w12540;
	assign w8857 = w45371 ^ w45246;
	assign w8615 = w8857 ^ w8791;
	assign w8626 = w8857 ^ w8798;
	assign w8575 = w45379 ^ w45246;
	assign w8870 = w8574 ^ w8575;
	assign w49603 = w45379 ^ w8615;
	assign w49579 = w45246 ^ w8655;
	assign w46908 = w49603 ^ w887;
	assign w30274 = w46908 ^ w46902;
	assign w30351 = w30268 ^ w30274;
	assign w30354 = w46903 ^ w30274;
	assign w46932 = w49579 ^ w863;
	assign w8638 = w8857 ^ w8845;
	assign w49595 = w45526 ^ w8626;
	assign w46916 = w49595 ^ w879;
	assign w27192 = w46916 ^ w46910;
	assign w27272 = w46911 ^ w27192;
	assign w27271 = w46916 ^ w27147;
	assign w27257 = w46916 & w27271;
	assign w16740 = w46932 ^ w46926;
	assign w16817 = w16734 ^ w16740;
	assign w16820 = w46927 ^ w16740;
	assign w12439 = w12435 ^ w12440;
	assign w12539 = w12438 ^ w12439;
	assign w49684 = ~w12539;
	assign w8856 = w45370 ^ w49684;
	assign w49596 = w8870 ^ w8856;
	assign w8567 = w12539 ^ w45371;
	assign w8873 = w8566 ^ w8567;
	assign w49580 = w8873 ^ w8845;
	assign w46915 = w49596 ^ w880;
	assign w27185 = w46915 ^ w46913;
	assign w27268 = w46915 ^ w27272;
	assign w27255 = w27272 & w27268;
	assign w46931 = w49580 ^ w864;
	assign w16733 = w46931 ^ w46929;
	assign w16814 = w16733 ^ w16822;
	assign w16735 = w46930 ^ w16733;
	assign w16810 = w16740 ^ w16735;
	assign w16811 = w46926 ^ w16735;
	assign w16813 = w46932 ^ w16814;
	assign w16808 = w46927 ^ w16735;
	assign w16750 = w46931 ^ w46930;
	assign w16815 = w16750 ^ w16817;
	assign w16823 = w46925 ^ w46931;
	assign w16818 = w16822 ^ w16750;
	assign w16801 = w16822 & w16811;
	assign w16709 = w16800 ^ w16801;
	assign w16737 = w16801 ^ w16735;
	assign w16807 = w16814 & w16818;
	assign w16739 = w16807 ^ w16736;
	assign w16806 = w16815 & w16813;
	assign w16804 = w16823 & w16808;
	assign w16738 = w16804 ^ w16734;
	assign w8636 = w8856 ^ w8841;
	assign w49589 = w49680 ^ w8636;
	assign w46922 = w49589 ^ w873;
	assign w11997 = w46917 ^ w46922;
	assign w16802 = w16817 & w16810;
	assign w16757 = w16800 ^ w16806;
	assign w16743 = w16739 ^ w16737;
	assign w16748 = w46925 ^ w16743;
	assign w16798 = w16757 ^ w16748;
	assign w8624 = w45378 ^ w12539;
	assign w49597 = w8623 ^ w8624;
	assign w46914 = w49597 ^ w881;
	assign w27187 = w46914 ^ w27185;
	assign w27263 = w46910 ^ w27187;
	assign w27260 = w46911 ^ w27187;
	assign w27262 = w27192 ^ w27187;
	assign w27202 = w46915 ^ w46914;
	assign w27276 = w46914 ^ w46912;
	assign w27162 = w46913 ^ w46914;
	assign w8614 = w8856 ^ w8853;
	assign w8612 = ~w8614;
	assign w16812 = w16733 ^ w16696;
	assign w16799 = w16821 & w16812;
	assign w44070 = w16799 ^ w16802;
	assign w16712 = w16738 ^ w44070;
	assign w16796 = w16712 ^ w16737;
	assign w16752 = w16800 ^ w44070;
	assign w16756 = w16709 ^ w16710;
	assign w16755 = w16756 ^ w16738;
	assign w16816 = w46931 ^ w16820;
	assign w16803 = w16820 & w16816;
	assign w16797 = w16803 ^ w16755;
	assign w16794 = w16798 & w16797;
	assign w16708 = w16803 ^ w16752;
	assign w16790 = w46931 ^ w16708;
	assign w16793 = w16794 ^ w16796;
	assign w11996 = w46919 ^ w11916;
	assign w45890 = ~w8794;
	assign w8633 = w45890 ^ w49682;
	assign w49591 = w8632 ^ w8633;
	assign w8639 = w45890 ^ w45370;
	assign w8637 = w8638 ^ w8639;
	assign w49588 = ~w8637;
	assign w46920 = w49591 ^ w875;
	assign w12000 = w46922 ^ w46920;
	assign w11912 = w46920 ^ w46918;
	assign w11871 = w11912 ^ w46919;
	assign w11985 = w11910 ^ w12000;
	assign w11976 = w12000 & w11985;
	assign w11872 = w11912 ^ w11910;
	assign w8616 = w45890 ^ w49698;
	assign w49602 = w8616 ^ w8617;
	assign w46909 = w49602 ^ w886;
	assign w27186 = w46911 ^ w46909;
	assign w27261 = w27186 ^ w27276;
	assign w27274 = w46912 ^ w46909;
	assign w27270 = w27274 ^ w27202;
	assign w27269 = w27186 ^ w27192;
	assign w27267 = w27202 ^ w27269;
	assign w27266 = w27185 ^ w27274;
	assign w27265 = w46916 ^ w27266;
	assign w27148 = w27188 ^ w27186;
	assign w27264 = w27185 ^ w27148;
	assign w27275 = w46909 ^ w46915;
	assign w27273 = w46909 ^ w46914;
	assign w27259 = w27266 & w27270;
	assign w27191 = w27259 ^ w27188;
	assign w27258 = w27267 & w27265;
	assign w27256 = w27275 & w27260;
	assign w27190 = w27256 ^ w27186;
	assign w27254 = w27269 & w27262;
	assign w27253 = w27274 & w27263;
	assign w27189 = w27253 ^ w27187;
	assign w27195 = w27191 ^ w27189;
	assign w27200 = w46909 ^ w27195;
	assign w27252 = w27276 & w27261;
	assign w27209 = w27252 ^ w27258;
	assign w27250 = w27209 ^ w27200;
	assign w27161 = w27252 ^ w27253;
	assign w27208 = w27161 ^ w27162;
	assign w27207 = w27208 ^ w27190;
	assign w27249 = w27255 ^ w27207;
	assign w27251 = w27273 & w27264;
	assign w27246 = w27250 & w27249;
	assign w44506 = w27251 ^ w27257;
	assign w27163 = w27195 ^ w44506;
	assign w27206 = w46911 ^ w27163;
	assign w27241 = w27246 ^ w27206;
	assign w27201 = w44506 ^ w27186;
	assign w27247 = w27209 ^ w27201;
	assign w44507 = w27251 ^ w27254;
	assign w27204 = w27252 ^ w44507;
	assign w27160 = w27255 ^ w27204;
	assign w27242 = w46915 ^ w27160;
	assign w27240 = w27241 & w27242;
	assign w27159 = w27240 ^ w27204;
	assign w27238 = w27246 ^ w27240;
	assign w27158 = w27240 ^ w27257;
	assign w27153 = w27158 ^ w27254;
	assign w27164 = w27190 ^ w44507;
	assign w27248 = w27164 ^ w27189;
	assign w27239 = w27240 ^ w27248;
	assign w27245 = w27246 ^ w27248;
	assign w27244 = w27247 & w27245;
	assign w27243 = w27244 ^ w27206;
	assign w27155 = w27244 ^ w27256;
	assign w27151 = w27155 ^ w27191;
	assign w27154 = w46909 ^ w27151;
	assign w27231 = w27153 ^ w27154;
	assign w27152 = w27244 ^ w27200;
	assign w27150 = w46911 ^ w27151;
	assign w27237 = w27248 & w27238;
	assign w27235 = w27237 ^ w27245;
	assign w27234 = w27243 & w27235;
	assign w27199 = w27234 ^ w27209;
	assign w27233 = w27199 ^ w27201;
	assign w27157 = w27234 ^ w27258;
	assign w27230 = w27199 ^ w27152;
	assign w27225 = w27239 & w46916;
	assign w27224 = w27230 & w27260;
	assign w27223 = w27233 & w27272;
	assign w27222 = w27243 & w27262;
	assign w27166 = w27222 ^ w27223;
	assign w27221 = w27231 & w27263;
	assign w27216 = w27239 & w27271;
	assign w27215 = w27230 & w27275;
	assign w27182 = w27224 ^ w27215;
	assign w27214 = w27233 & w27268;
	assign w27184 = w27222 ^ w27214;
	assign w27213 = w27243 & w27269;
	assign w27212 = w27231 & w27274;
	assign w44509 = w27223 ^ w27224;
	assign w44511 = w27237 ^ w27255;
	assign w27229 = w44511 ^ w27207;
	assign w27227 = w27229 & w27266;
	assign w44510 = w27225 ^ w27227;
	assign w27218 = w27229 & w27270;
	assign w27196 = w46915 ^ w44511;
	assign w27236 = w27196 ^ w27159;
	assign w27149 = w27196 ^ w27157;
	assign w27156 = w27186 ^ w27149;
	assign w27232 = w27153 ^ w27156;
	assign w27228 = w27149 ^ w27150;
	assign w27226 = w27236 & w27265;
	assign w27220 = w27228 & w27261;
	assign w27205 = w27220 ^ w44509;
	assign w27181 = w27220 ^ w27223;
	assign w27178 = ~w27181;
	assign w27177 = w27220 ^ w27221;
	assign w27171 = w27216 ^ w27205;
	assign w27168 = ~w27171;
	assign w27165 = w27221 ^ w27205;
	assign w27219 = w27232 & w27264;
	assign w27197 = w27215 ^ w27219;
	assign w27175 = ~w27197;
	assign w27174 = w27175 ^ w27213;
	assign w27170 = w27174 ^ w44510;
	assign w27173 = w27212 ^ w27170;
	assign w27217 = w27236 & w27267;
	assign w27211 = w27228 & w27276;
	assign w27210 = w27232 & w27273;
	assign w27176 = w27221 ^ w27210;
	assign w27172 = ~w27176;
	assign w27277 = w27172 ^ w27173;
	assign w44508 = w27211 ^ w27212;
	assign w27193 = w27217 ^ w44508;
	assign w27169 = w27193 ^ w27170;
	assign w49909 = w27168 ^ w27169;
	assign w27194 = w27218 ^ w27193;
	assign w49912 = w27194 ^ w27165;
	assign w27198 = w27226 ^ w27194;
	assign w27167 = w27225 ^ w27198;
	assign w49910 = w27166 ^ w27167;
	assign w27203 = w27227 ^ w27198;
	assign w27278 = w27203 ^ w27177;
	assign w49911 = w44509 ^ w27203;
	assign w27180 = w27184 ^ w44508;
	assign w27183 = w44510 ^ w27180;
	assign w27280 = w27182 ^ w27183;
	assign w27179 = w27175 ^ w27180;
	assign w27279 = w27178 ^ w27179;
	assign w11995 = w46924 ^ w11871;
	assign w11981 = w46924 & w11995;
	assign w8635 = w45890 ^ w49681;
	assign w49590 = w8634 ^ w8635;
	assign w46921 = w49590 ^ w874;
	assign w11886 = w46921 ^ w46922;
	assign w46923 = w49588 ^ w872;
	assign w11999 = w46917 ^ w46923;
	assign w11992 = w46923 ^ w11996;
	assign w11909 = w46923 ^ w46921;
	assign w11911 = w46922 ^ w11909;
	assign w11986 = w11916 ^ w11911;
	assign w11978 = w11993 & w11986;
	assign w11988 = w11909 ^ w11872;
	assign w11975 = w11997 & w11988;
	assign w11926 = w46923 ^ w46922;
	assign w11991 = w11926 ^ w11993;
	assign w11987 = w46918 ^ w11911;
	assign w11984 = w46919 ^ w11911;
	assign w11980 = w11999 & w11984;
	assign w11914 = w11980 ^ w11910;
	assign w43869 = w11975 ^ w11978;
	assign w11888 = w11914 ^ w43869;
	assign w11928 = w11976 ^ w43869;
	assign w43872 = w11975 ^ w11981;
	assign w11925 = w43872 ^ w11910;
	assign w11998 = w46920 ^ w46917;
	assign w11994 = w11998 ^ w11926;
	assign w11977 = w11998 & w11987;
	assign w11913 = w11977 ^ w11911;
	assign w11972 = w11888 ^ w11913;
	assign w11885 = w11976 ^ w11977;
	assign w11932 = w11885 ^ w11886;
	assign w11990 = w11909 ^ w11998;
	assign w11983 = w11990 & w11994;
	assign w11989 = w46924 ^ w11990;
	assign w11982 = w11991 & w11989;
	assign w11933 = w11976 ^ w11982;
	assign w11971 = w11933 ^ w11925;
	assign w11931 = w11932 ^ w11914;
	assign w11915 = w11983 ^ w11912;
	assign w11919 = w11915 ^ w11913;
	assign w11887 = w11919 ^ w43872;
	assign w11924 = w46917 ^ w11919;
	assign w11930 = w46919 ^ w11887;
	assign w11974 = w11933 ^ w11924;
	assign w8941 = w49911 ^ w49910;
	assign w45606 = ~w27278;
	assign w45607 = ~w27279;
	assign w45608 = ~w27280;
	assign w45613 = ~w27277;
	assign w9089 = w45606 ^ w45613;
	assign w11979 = w11996 & w11992;
	assign w11884 = w11979 ^ w11928;
	assign w11966 = w46923 ^ w11884;
	assign w11973 = w11979 ^ w11931;
	assign w11970 = w11974 & w11973;
	assign w11965 = w11970 ^ w11930;
	assign w11964 = w11965 & w11966;
	assign w11883 = w11964 ^ w11928;
	assign w11882 = w11964 ^ w11981;
	assign w11877 = w11882 ^ w11978;
	assign w11962 = w11970 ^ w11964;
	assign w11961 = w11972 & w11962;
	assign w11963 = w11964 ^ w11972;
	assign w11949 = w11963 & w46924;
	assign w11940 = w11963 & w11995;
	assign w43871 = w11961 ^ w11979;
	assign w11920 = w46923 ^ w43871;
	assign w11960 = w11920 ^ w11883;
	assign w11941 = w11960 & w11991;
	assign w11950 = w11960 & w11989;
	assign w11953 = w43871 ^ w11931;
	assign w11942 = w11953 & w11994;
	assign w11951 = w11953 & w11990;
	assign w43874 = w11949 ^ w11951;
	assign w11969 = w11970 ^ w11972;
	assign w11968 = w11971 & w11969;
	assign w11879 = w11968 ^ w11980;
	assign w11875 = w11879 ^ w11915;
	assign w11878 = w46917 ^ w11875;
	assign w11967 = w11968 ^ w11930;
	assign w11946 = w11967 & w11986;
	assign w11955 = w11877 ^ w11878;
	assign w11936 = w11955 & w11998;
	assign w11945 = w11955 & w11987;
	assign w11959 = w11961 ^ w11969;
	assign w11958 = w11967 & w11959;
	assign w11881 = w11958 ^ w11982;
	assign w11873 = w11920 ^ w11881;
	assign w11880 = w11910 ^ w11873;
	assign w11923 = w11958 ^ w11933;
	assign w11957 = w11923 ^ w11925;
	assign w11947 = w11957 & w11996;
	assign w11938 = w11957 & w11992;
	assign w11908 = w11946 ^ w11938;
	assign w11956 = w11877 ^ w11880;
	assign w11943 = w11956 & w11988;
	assign w11876 = w11968 ^ w11924;
	assign w11937 = w11967 & w11993;
	assign w11954 = w11923 ^ w11876;
	assign w11948 = w11954 & w11984;
	assign w11939 = w11954 & w11999;
	assign w11906 = w11948 ^ w11939;
	assign w11921 = w11939 ^ w11943;
	assign w11899 = ~w11921;
	assign w11898 = w11899 ^ w11937;
	assign w11894 = w11898 ^ w43874;
	assign w11897 = w11936 ^ w11894;
	assign w11874 = w46919 ^ w11875;
	assign w11952 = w11873 ^ w11874;
	assign w11944 = w11952 & w11985;
	assign w11935 = w11952 & w12000;
	assign w11905 = w11944 ^ w11947;
	assign w11902 = ~w11905;
	assign w11901 = w11944 ^ w11945;
	assign w43870 = w11935 ^ w11936;
	assign w11917 = w11941 ^ w43870;
	assign w11893 = w11917 ^ w11894;
	assign w43873 = w11947 ^ w11948;
	assign w11929 = w11944 ^ w43873;
	assign w11895 = w11940 ^ w11929;
	assign w11892 = ~w11895;
	assign w49848 = w11892 ^ w11893;
	assign w8931 = w49844 ^ w49848;
	assign w11889 = w11945 ^ w11929;
	assign w11934 = w11956 & w11997;
	assign w11900 = w11945 ^ w11934;
	assign w11896 = ~w11900;
	assign w11904 = w11908 ^ w43870;
	assign w11903 = w11899 ^ w11904;
	assign w12003 = w11902 ^ w11903;
	assign w11907 = w43874 ^ w11904;
	assign w12004 = w11906 ^ w11907;
	assign w45240 = ~w12003;
	assign w45241 = ~w12004;
	assign w12001 = w11896 ^ w11897;
	assign w49851 = ~w12001;
	assign w9192 = w45617 ^ w49851;
	assign w11918 = w11942 ^ w11917;
	assign w11922 = w11950 ^ w11918;
	assign w11891 = w11949 ^ w11922;
	assign w49853 = w11918 ^ w11889;
	assign w9140 = w49847 ^ w49853;
	assign w8930 = w9140 ^ w49845;
	assign w11927 = w11951 ^ w11922;
	assign w49850 = w43873 ^ w11927;
	assign w9195 = w49846 ^ w49850;
	assign w9209 = w8930 ^ w8931;
	assign w12002 = w11927 ^ w11901;
	assign w49852 = ~w12002;
	assign w9190 = w45610 ^ w49852;
	assign w11890 = w11946 ^ w11947;
	assign w49849 = w11890 ^ w11891;
	assign w9204 = w49845 ^ w49849;
	assign w9086 = ~w9204;
	assign w16695 = w16736 ^ w46927;
	assign w16819 = w46932 ^ w16695;
	assign w16805 = w46932 & w16819;
	assign w44073 = w16799 ^ w16805;
	assign w16749 = w44073 ^ w16734;
	assign w16795 = w16757 ^ w16749;
	assign w16792 = w16795 & w16793;
	assign w16703 = w16792 ^ w16804;
	assign w16699 = w16703 ^ w16739;
	assign w16698 = w46927 ^ w16699;
	assign w16700 = w16792 ^ w16748;
	assign w16711 = w16743 ^ w44073;
	assign w16754 = w46927 ^ w16711;
	assign w16791 = w16792 ^ w16754;
	assign w16789 = w16794 ^ w16754;
	assign w16770 = w16791 & w16810;
	assign w16761 = w16791 & w16817;
	assign w16702 = w46925 ^ w16699;
	assign w16788 = w16789 & w16790;
	assign w16786 = w16794 ^ w16788;
	assign w16785 = w16796 & w16786;
	assign w16783 = w16785 ^ w16793;
	assign w16782 = w16791 & w16783;
	assign w16787 = w16788 ^ w16796;
	assign w16773 = w16787 & w46932;
	assign w16764 = w16787 & w16819;
	assign w16706 = w16788 ^ w16805;
	assign w16701 = w16706 ^ w16802;
	assign w16779 = w16701 ^ w16702;
	assign w16769 = w16779 & w16811;
	assign w16760 = w16779 & w16822;
	assign w16705 = w16782 ^ w16806;
	assign w16707 = w16788 ^ w16752;
	assign w16747 = w16782 ^ w16757;
	assign w16778 = w16747 ^ w16700;
	assign w16772 = w16778 & w16808;
	assign w16781 = w16747 ^ w16749;
	assign w16762 = w16781 & w16816;
	assign w16771 = w16781 & w16820;
	assign w16763 = w16778 & w16823;
	assign w16730 = w16772 ^ w16763;
	assign w16732 = w16770 ^ w16762;
	assign w16714 = w16770 ^ w16771;
	assign w44072 = w16785 ^ w16803;
	assign w16777 = w44072 ^ w16755;
	assign w16775 = w16777 & w16814;
	assign w16766 = w16777 & w16818;
	assign w16744 = w46931 ^ w44072;
	assign w16697 = w16744 ^ w16705;
	assign w16776 = w16697 ^ w16698;
	assign w16768 = w16776 & w16809;
	assign w16729 = w16768 ^ w16771;
	assign w16726 = ~w16729;
	assign w16725 = w16768 ^ w16769;
	assign w16784 = w16744 ^ w16707;
	assign w16765 = w16784 & w16815;
	assign w16774 = w16784 & w16813;
	assign w44074 = w16771 ^ w16772;
	assign w16753 = w16768 ^ w44074;
	assign w16719 = w16764 ^ w16753;
	assign w16716 = ~w16719;
	assign w44075 = w16773 ^ w16775;
	assign w16704 = w16734 ^ w16697;
	assign w16759 = w16776 & w16824;
	assign w44071 = w16759 ^ w16760;
	assign w16728 = w16732 ^ w44071;
	assign w16731 = w44075 ^ w16728;
	assign w16828 = w16730 ^ w16731;
	assign w45350 = ~w16828;
	assign w16741 = w16765 ^ w44071;
	assign w16742 = w16766 ^ w16741;
	assign w16746 = w16774 ^ w16742;
	assign w16715 = w16773 ^ w16746;
	assign w49865 = w16714 ^ w16715;
	assign w16751 = w16775 ^ w16746;
	assign w49866 = w44074 ^ w16751;
	assign w16826 = w16751 ^ w16725;
	assign w45356 = ~w16826;
	assign w9155 = w45356 ^ w45523;
	assign w16780 = w16701 ^ w16704;
	assign w16767 = w16780 & w16812;
	assign w16745 = w16763 ^ w16767;
	assign w16758 = w16780 & w16821;
	assign w16724 = w16769 ^ w16758;
	assign w16720 = ~w16724;
	assign w16723 = ~w16745;
	assign w16727 = w16723 ^ w16728;
	assign w16827 = w16726 ^ w16727;
	assign w16722 = w16723 ^ w16761;
	assign w16718 = w16722 ^ w44075;
	assign w16717 = w16741 ^ w16718;
	assign w49864 = w16716 ^ w16717;
	assign w16721 = w16760 ^ w16718;
	assign w16825 = w16720 ^ w16721;
	assign w45355 = ~w16825;
	assign w45357 = ~w16827;
	assign w16713 = w16769 ^ w16753;
	assign w49867 = w16742 ^ w16713;
	assign w9146 = w49867 ^ w49880;
	assign w9028 = w49867 ^ w45356;
	assign w8893 = ~w9146;
	assign w8894 = w8893 ^ w49877;
	assign w8891 = w8893 ^ w45525;
	assign w8897 = w9146 ^ w49878;
	assign w24195 = w24090 ^ w24091;
	assign w45522 = ~w24195;
	assign w9047 = w45522 ^ w45355;
	assign w45932 = ~w8451;
	assign w8283 = w45932 ^ w45403;
	assign w49321 = w8283 ^ w8284;
	assign w8370 = w45932 ^ w49455;
	assign w49342 = w8369 ^ w8370;
	assign w8246 = w45932 ^ w49457;
	assign w8519 = w8246 ^ w8247;
	assign w49341 = w8519 ^ w8516;
	assign w47097 = w49341 ^ w1846;
	assign w30669 = w47099 ^ w47097;
	assign w30671 = w47098 ^ w30669;
	assign w30747 = w47094 ^ w30671;
	assign w30744 = w47095 ^ w30671;
	assign w30746 = w30676 ^ w30671;
	assign w30646 = w47097 ^ w47098;
	assign w30740 = w30759 & w30744;
	assign w30674 = w30740 ^ w30670;
	assign w30738 = w30753 & w30746;
	assign w47117 = w49321 ^ w1826;
	assign w18028 = w47120 ^ w47117;
	assign w18020 = w17939 ^ w18028;
	assign w17940 = w47119 ^ w47117;
	assign w18023 = w17940 ^ w17946;
	assign w18008 = w18023 & w18016;
	assign w18007 = w18028 & w18017;
	assign w17943 = w18007 ^ w17941;
	assign w17902 = w17942 ^ w17940;
	assign w18015 = w17940 ^ w18030;
	assign w18006 = w18030 & w18015;
	assign w17915 = w18006 ^ w18007;
	assign w17962 = w17915 ^ w17916;
	assign w18021 = w17956 ^ w18023;
	assign w47096 = w49342 ^ w1847;
	assign w30672 = w47096 ^ w47094;
	assign w30758 = w47096 ^ w47093;
	assign w30754 = w30758 ^ w30686;
	assign w30750 = w30669 ^ w30758;
	assign w30749 = w47100 ^ w30750;
	assign w30760 = w47098 ^ w47096;
	assign w30745 = w30670 ^ w30760;
	assign w30632 = w30672 ^ w30670;
	assign w30748 = w30669 ^ w30632;
	assign w30631 = w30672 ^ w47095;
	assign w30755 = w47100 ^ w30631;
	assign w30743 = w30750 & w30754;
	assign w30675 = w30743 ^ w30672;
	assign w30742 = w30751 & w30749;
	assign w30741 = w47100 & w30755;
	assign w30737 = w30758 & w30747;
	assign w30673 = w30737 ^ w30671;
	assign w30679 = w30675 ^ w30673;
	assign w30684 = w47093 ^ w30679;
	assign w30736 = w30760 & w30745;
	assign w30693 = w30736 ^ w30742;
	assign w30734 = w30693 ^ w30684;
	assign w30645 = w30736 ^ w30737;
	assign w30692 = w30645 ^ w30646;
	assign w30691 = w30692 ^ w30674;
	assign w30733 = w30739 ^ w30691;
	assign w30735 = w30757 & w30748;
	assign w30730 = w30734 & w30733;
	assign w18018 = w17939 ^ w17902;
	assign w44654 = w30735 ^ w30741;
	assign w30647 = w30679 ^ w44654;
	assign w30690 = w47095 ^ w30647;
	assign w30725 = w30730 ^ w30690;
	assign w30685 = w44654 ^ w30670;
	assign w30731 = w30693 ^ w30685;
	assign w44655 = w30735 ^ w30738;
	assign w30688 = w30736 ^ w44655;
	assign w30644 = w30739 ^ w30688;
	assign w30726 = w47099 ^ w30644;
	assign w30724 = w30725 & w30726;
	assign w30643 = w30724 ^ w30688;
	assign w30642 = w30724 ^ w30741;
	assign w30637 = w30642 ^ w30738;
	assign w30722 = w30730 ^ w30724;
	assign w30648 = w30674 ^ w44655;
	assign w30732 = w30648 ^ w30673;
	assign w30723 = w30724 ^ w30732;
	assign w30729 = w30730 ^ w30732;
	assign w30728 = w30731 & w30729;
	assign w30727 = w30728 ^ w30690;
	assign w30639 = w30728 ^ w30740;
	assign w30635 = w30639 ^ w30675;
	assign w30638 = w47093 ^ w30635;
	assign w30715 = w30637 ^ w30638;
	assign w30636 = w30728 ^ w30684;
	assign w30634 = w47095 ^ w30635;
	assign w30721 = w30732 & w30722;
	assign w30719 = w30721 ^ w30729;
	assign w30718 = w30727 & w30719;
	assign w30683 = w30718 ^ w30693;
	assign w30717 = w30683 ^ w30685;
	assign w30641 = w30718 ^ w30742;
	assign w30714 = w30683 ^ w30636;
	assign w30709 = w30723 & w47100;
	assign w30708 = w30714 & w30744;
	assign w30707 = w30717 & w30756;
	assign w30706 = w30727 & w30746;
	assign w30650 = w30706 ^ w30707;
	assign w30705 = w30715 & w30747;
	assign w30700 = w30723 & w30755;
	assign w30699 = w30714 & w30759;
	assign w30666 = w30708 ^ w30699;
	assign w30698 = w30717 & w30752;
	assign w30668 = w30706 ^ w30698;
	assign w30697 = w30727 & w30753;
	assign w30696 = w30715 & w30758;
	assign w44657 = w30707 ^ w30708;
	assign w44659 = w30721 ^ w30739;
	assign w30713 = w44659 ^ w30691;
	assign w30711 = w30713 & w30750;
	assign w44658 = w30709 ^ w30711;
	assign w30702 = w30713 & w30754;
	assign w30680 = w47099 ^ w44659;
	assign w30720 = w30680 ^ w30643;
	assign w30633 = w30680 ^ w30641;
	assign w30640 = w30670 ^ w30633;
	assign w30716 = w30637 ^ w30640;
	assign w30712 = w30633 ^ w30634;
	assign w30710 = w30720 & w30749;
	assign w30704 = w30712 & w30745;
	assign w30689 = w30704 ^ w44657;
	assign w30665 = w30704 ^ w30707;
	assign w30662 = ~w30665;
	assign w30661 = w30704 ^ w30705;
	assign w30655 = w30700 ^ w30689;
	assign w30652 = ~w30655;
	assign w30649 = w30705 ^ w30689;
	assign w30703 = w30716 & w30748;
	assign w30681 = w30699 ^ w30703;
	assign w30659 = ~w30681;
	assign w30658 = w30659 ^ w30697;
	assign w30654 = w30658 ^ w44658;
	assign w30657 = w30696 ^ w30654;
	assign w30701 = w30720 & w30751;
	assign w30695 = w30712 & w30760;
	assign w30694 = w30716 & w30757;
	assign w30660 = w30705 ^ w30694;
	assign w30656 = ~w30660;
	assign w30761 = w30656 ^ w30657;
	assign w44656 = w30695 ^ w30696;
	assign w30677 = w30701 ^ w44656;
	assign w30653 = w30677 ^ w30654;
	assign w49658 = w30652 ^ w30653;
	assign w30678 = w30702 ^ w30677;
	assign w49662 = w30678 ^ w30649;
	assign w8803 = w49646 ^ w49662;
	assign w30682 = w30710 ^ w30678;
	assign w30651 = w30709 ^ w30682;
	assign w49659 = w30650 ^ w30651;
	assign w30687 = w30711 ^ w30682;
	assign w30762 = w30687 ^ w30661;
	assign w49661 = ~w30762;
	assign w8840 = w45528 ^ w49661;
	assign w8788 = w8836 ^ w8803;
	assign w8850 = w49655 ^ w49659;
	assign w49526 = w8865 ^ w8850;
	assign w8545 = w8803 ^ w49644;
	assign w8546 = w49659 ^ w49649;
	assign w8882 = w8545 ^ w8546;
	assign w8647 = w8840 ^ w45388;
	assign w8730 = w8731 ^ w49659;
	assign w49534 = w8729 ^ w8730;
	assign w8722 = w8846 ^ w30762;
	assign w8699 = ~w8803;
	assign w49537 = w8722 ^ w8723;
	assign w8698 = w8699 ^ w49648;
	assign w8738 = w8848 ^ w8840;
	assign w49529 = w45389 ^ w8738;
	assign w8709 = w8840 ^ w8796;
	assign w49546 = w49657 ^ w8709;
	assign w46965 = w49546 ^ w958;
	assign w46977 = w49534 ^ w946;
	assign w8838 = w49643 ^ w49658;
	assign w8732 = w8838 ^ w8837;
	assign w49533 = w49647 ^ w8732;
	assign w8700 = ~w8838;
	assign w8697 = w8850 ^ w8700;
	assign w49518 = w8697 ^ w8698;
	assign w8769 = w8700 ^ w45247;
	assign w49525 = w8769 ^ w8770;
	assign w46986 = w49525 ^ w937;
	assign w8715 = w8851 ^ w8850;
	assign w8713 = ~w8715;
	assign w8628 = w30762 ^ w49652;
	assign w46985 = w49526 ^ w938;
	assign w33326 = w46985 ^ w46986;
	assign w46993 = w49518 ^ w930;
	assign w46978 = w49533 ^ w945;
	assign w16978 = w46977 ^ w46978;
	assign w8795 = w49657 ^ w49662;
	assign w8719 = w8836 ^ w8795;
	assign w49539 = w45383 ^ w8719;
	assign w8737 = w8846 ^ w8795;
	assign w49530 = w49646 ^ w8737;
	assign w46981 = w49530 ^ w942;
	assign w33437 = w46981 ^ w46986;
	assign w46974 = w49537 ^ w949;
	assign w46982 = w49529 ^ w941;
	assign w49660 = w44657 ^ w30687;
	assign w8847 = w49656 ^ w49660;
	assign w8712 = w8848 ^ w8847;
	assign w49544 = w45527 ^ w8712;
	assign w49519 = w8882 ^ w8847;
	assign w46992 = w49519 ^ w931;
	assign w46967 = w49544 ^ w956;
	assign w30402 = w46967 ^ w46965;
	assign w8740 = w8742 ^ w8847;
	assign w8582 = w8797 ^ w49660;
	assign w8867 = w8582 ^ w8583;
	assign w49535 = w8867 ^ w8851;
	assign w46976 = w49535 ^ w947;
	assign w17004 = w46976 ^ w46974;
	assign w17092 = w46978 ^ w46976;
	assign w8665 = w49660 ^ w12403;
	assign w30664 = w30668 ^ w44656;
	assign w30667 = w44658 ^ w30664;
	assign w30764 = w30666 ^ w30667;
	assign w30663 = w30659 ^ w30664;
	assign w30763 = w30662 ^ w30663;
	assign w18027 = w47117 ^ w47122;
	assign w18005 = w18027 & w18018;
	assign w44120 = w18005 ^ w18008;
	assign w17958 = w18006 ^ w44120;
	assign w17914 = w18009 ^ w17958;
	assign w17996 = w47123 ^ w17914;
	assign w44123 = w18005 ^ w18011;
	assign w17955 = w44123 ^ w17940;
	assign w18029 = w47117 ^ w47123;
	assign w18010 = w18029 & w18014;
	assign w46972 = w49539 ^ w951;
	assign w17944 = w18010 ^ w17940;
	assign w17918 = w17944 ^ w44120;
	assign w18002 = w17918 ^ w17943;
	assign w17961 = w17962 ^ w17944;
	assign w18003 = w18009 ^ w17961;
	assign w18024 = w18028 ^ w17956;
	assign w18013 = w18020 & w18024;
	assign w17945 = w18013 ^ w17942;
	assign w17949 = w17945 ^ w17943;
	assign w17917 = w17949 ^ w44123;
	assign w17960 = w47119 ^ w17917;
	assign w17954 = w47117 ^ w17949;
	assign w18019 = w47124 ^ w18020;
	assign w18012 = w18021 & w18019;
	assign w17963 = w18006 ^ w18012;
	assign w18004 = w17963 ^ w17954;
	assign w18000 = w18004 & w18003;
	assign w17999 = w18000 ^ w18002;
	assign w17995 = w18000 ^ w17960;
	assign w17994 = w17995 & w17996;
	assign w17913 = w17994 ^ w17958;
	assign w17912 = w17994 ^ w18011;
	assign w17907 = w17912 ^ w18008;
	assign w17993 = w17994 ^ w18002;
	assign w17970 = w17993 & w18025;
	assign w17979 = w17993 & w47124;
	assign w17992 = w18000 ^ w17994;
	assign w17991 = w18002 & w17992;
	assign w44122 = w17991 ^ w18009;
	assign w17983 = w44122 ^ w17961;
	assign w17981 = w17983 & w18020;
	assign w17972 = w17983 & w18024;
	assign w17950 = w47123 ^ w44122;
	assign w17990 = w17950 ^ w17913;
	assign w17971 = w17990 & w18021;
	assign w44125 = w17979 ^ w17981;
	assign w17980 = w17990 & w18019;
	assign w17989 = w17991 ^ w17999;
	assign w18001 = w17963 ^ w17955;
	assign w17998 = w18001 & w17999;
	assign w17906 = w17998 ^ w17954;
	assign w17909 = w17998 ^ w18010;
	assign w17905 = w17909 ^ w17945;
	assign w17904 = w47119 ^ w17905;
	assign w17908 = w47117 ^ w17905;
	assign w17997 = w17998 ^ w17960;
	assign w17988 = w17997 & w17989;
	assign w17976 = w17997 & w18016;
	assign w17911 = w17988 ^ w18012;
	assign w17967 = w17997 & w18023;
	assign w17953 = w17988 ^ w17963;
	assign w17984 = w17953 ^ w17906;
	assign w17969 = w17984 & w18029;
	assign w17987 = w17953 ^ w17955;
	assign w17977 = w17987 & w18026;
	assign w17920 = w17976 ^ w17977;
	assign w17978 = w17984 & w18014;
	assign w17936 = w17978 ^ w17969;
	assign w17968 = w17987 & w18022;
	assign w17938 = w17976 ^ w17968;
	assign w44124 = w17977 ^ w17978;
	assign w17903 = w17950 ^ w17911;
	assign w17910 = w17940 ^ w17903;
	assign w17982 = w17903 ^ w17904;
	assign w17965 = w17982 & w18030;
	assign w17986 = w17907 ^ w17910;
	assign w17974 = w17982 & w18015;
	assign w17959 = w17974 ^ w44124;
	assign w17925 = w17970 ^ w17959;
	assign w17922 = ~w17925;
	assign w17935 = w17974 ^ w17977;
	assign w17973 = w17986 & w18018;
	assign w17951 = w17969 ^ w17973;
	assign w17929 = ~w17951;
	assign w17928 = w17929 ^ w17967;
	assign w17985 = w17907 ^ w17908;
	assign w17975 = w17985 & w18017;
	assign w17931 = w17974 ^ w17975;
	assign w17919 = w17975 ^ w17959;
	assign w17966 = w17985 & w18028;
	assign w44121 = w17965 ^ w17966;
	assign w17947 = w17971 ^ w44121;
	assign w17934 = w17938 ^ w44121;
	assign w17937 = w44125 ^ w17934;
	assign w17933 = w17929 ^ w17934;
	assign w18034 = w17936 ^ w17937;
	assign w17964 = w17986 & w18027;
	assign w17930 = w17975 ^ w17964;
	assign w17926 = ~w17930;
	assign w17948 = w17972 ^ w17947;
	assign w49703 = w17948 ^ w17919;
	assign w8801 = w49703 ^ w49715;
	assign w8787 = w8801 ^ w49706;
	assign w8600 = w8839 ^ w8801;
	assign w49611 = w45776 ^ w8600;
	assign w46900 = w49611 ^ w1851;
	assign w8790 = w49703 ^ w49707;
	assign w8755 = w8790 ^ w49715;
	assign w49634 = w8755 ^ w8756;
	assign w8743 = w8812 ^ w8790;
	assign w49642 = w49711 ^ w8743;
	assign w46869 = w49642 ^ w1882;
	assign w8779 = w8839 ^ w8790;
	assign w46877 = w49634 ^ w1874;
	assign w45387 = ~w18034;
	assign w8852 = w45387 ^ w45776;
	assign w8555 = w8801 ^ w45387;
	assign w8878 = w8555 ^ w8556;
	assign w49612 = w8878 ^ w8819;
	assign w8754 = w8852 ^ w8789;
	assign w49635 = w45375 ^ w8754;
	assign w8777 = w8852 ^ w8819;
	assign w49619 = w45387 ^ w8779;
	assign w46892 = w49619 ^ w1859;
	assign w46876 = w49635 ^ w1875;
	assign w46899 = w49612 ^ w1852;
	assign w8764 = w8852 ^ w8804;
	assign w49627 = w45367 ^ w8764;
	assign w46884 = w49627 ^ w1867;
	assign w17952 = w17980 ^ w17948;
	assign w17957 = w17981 ^ w17952;
	assign w18032 = w17957 ^ w17931;
	assign w8781 = w49707 ^ w18032;
	assign w49702 = ~w18032;
	assign w8854 = w49702 ^ w45774;
	assign w8765 = w8854 ^ w8789;
	assign w8757 = w8854 ^ w8814;
	assign w49633 = w45373 ^ w8757;
	assign w17921 = w17979 ^ w17952;
	assign w49700 = w17920 ^ w17921;
	assign w8815 = w49700 ^ w49713;
	assign w8786 = w8815 ^ w8806;
	assign w49630 = w8883 ^ w8815;
	assign w8744 = w8854 ^ w45372;
	assign w49641 = w8744 ^ w8745;
	assign w46870 = w49641 ^ w1881;
	assign w30140 = w46876 ^ w46870;
	assign w49615 = w8786 ^ w8787;
	assign w46896 = w49615 ^ w1855;
	assign w49701 = w44124 ^ w17957;
	assign w8855 = w49701 ^ w49706;
	assign w49639 = w8861 ^ w8855;
	assign w8760 = w8855 ^ w8809;
	assign w46872 = w49639 ^ w1879;
	assign w30136 = w46872 ^ w46870;
	assign w30222 = w46872 ^ w46869;
	assign w8595 = ~w49701;
	assign w8594 = w49705 ^ w8595;
	assign w8784 = w49714 ^ w8595;
	assign w49616 = w8783 ^ w8784;
	assign w46895 = w49616 ^ w1856;
	assign w46878 = w49633 ^ w1873;
	assign w46881 = w49630 ^ w1870;
	assign w49631 = w8760 ^ w8761;
	assign w46880 = w49631 ^ w1871;
	assign w16468 = w46880 ^ w46878;
	assign w49626 = w49703 ^ w8765;
	assign w46885 = w49626 ^ w1866;
	assign w16472 = w46884 ^ w46878;
	assign w17932 = ~w17935;
	assign w18033 = w17932 ^ w17933;
	assign w45386 = ~w18033;
	assign w8844 = w45386 ^ w45775;
	assign w8598 = w8807 ^ w45386;
	assign w49613 = w8598 ^ w8599;
	assign w8753 = ~w8844;
	assign w8751 = w8753 ^ w8839;
	assign w46898 = w49613 ^ w1853;
	assign w16616 = w46899 ^ w46898;
	assign w8775 = w8844 ^ w8807;
	assign w49628 = w8884 ^ w8844;
	assign w46883 = w49628 ^ w1868;
	assign w16465 = w46883 ^ w46881;
	assign w16555 = w46877 ^ w46883;
	assign w16690 = w46898 ^ w46896;
	assign w45702 = ~w30764;
	assign w8859 = w45383 ^ w45702;
	assign w49515 = w45702 ^ w8788;
	assign w8588 = w8795 ^ w45702;
	assign w8864 = w8588 ^ w8589;
	assign w8611 = w8859 ^ w8796;
	assign w49523 = w45529 ^ w8611;
	assign w8727 = w8859 ^ w8837;
	assign w8736 = w8859 ^ w8797;
	assign w49531 = w45248 ^ w8736;
	assign w46988 = w49523 ^ w935;
	assign w33356 = w46988 ^ w46982;
	assign w46980 = w49531 ^ w943;
	assign w46996 = w49515 ^ w927;
	assign w17008 = w46980 ^ w46974;
	assign w49540 = w8864 ^ w8837;
	assign w46971 = w49540 ^ w952;
	assign w30491 = w46965 ^ w46971;
	assign w45708 = ~w30761;
	assign w8724 = w8848 ^ w45708;
	assign w49536 = w8724 ^ w8725;
	assign w8648 = w45708 ^ w12404;
	assign w8646 = w8647 ^ w8648;
	assign w49521 = ~w8646;
	assign w46975 = w49536 ^ w948;
	assign w16963 = w17004 ^ w46975;
	assign w17087 = w46980 ^ w16963;
	assign w17073 = w46980 & w17087;
	assign w17088 = w46975 ^ w17008;
	assign w46990 = w49521 ^ w933;
	assign w17138 = w46992 ^ w46990;
	assign w17142 = w46996 ^ w46990;
	assign w8843 = w45527 ^ w45708;
	assign w8666 = w8843 ^ w49645;
	assign w8664 = ~w8666;
	assign w49520 = w8664 ^ w8665;
	assign w8710 = w8846 ^ w8843;
	assign w8739 = w8851 ^ w8843;
	assign w49528 = w45388 ^ w8739;
	assign w49545 = w45528 ^ w8710;
	assign w46966 = w49545 ^ w957;
	assign w30408 = w46972 ^ w46966;
	assign w30485 = w30402 ^ w30408;
	assign w30488 = w46967 ^ w30408;
	assign w30484 = w46971 ^ w30488;
	assign w30471 = w30488 & w30484;
	assign w46983 = w49528 ^ w940;
	assign w33350 = w46983 ^ w46981;
	assign w33433 = w33350 ^ w33356;
	assign w33436 = w46983 ^ w33356;
	assign w46991 = w49520 ^ w932;
	assign w17222 = w46991 ^ w17142;
	assign w17097 = w17138 ^ w46991;
	assign w17221 = w46996 ^ w17097;
	assign w17207 = w46996 & w17221;
	assign w45709 = ~w30763;
	assign w8858 = w45382 ^ w45709;
	assign w8728 = w8699 ^ w45709;
	assign w8726 = w8727 ^ w8728;
	assign w8717 = w45709 ^ w24331;
	assign w49516 = ~w8726;
	assign w49541 = w8716 ^ w8717;
	assign w8711 = w8858 ^ w8835;
	assign w49517 = w49658 ^ w8711;
	assign w46994 = w49517 ^ w929;
	assign w17226 = w46994 ^ w46992;
	assign w17112 = w46993 ^ w46994;
	assign w46995 = w49516 ^ w928;
	assign w17135 = w46995 ^ w46993;
	assign w17218 = w46995 ^ w17222;
	assign w17152 = w46995 ^ w46994;
	assign w17205 = w17222 & w17218;
	assign w46970 = w49541 ^ w953;
	assign w30418 = w46971 ^ w46970;
	assign w30483 = w30418 ^ w30485;
	assign w30489 = w46965 ^ w46970;
	assign w8734 = w8858 ^ w8836;
	assign w17137 = w46994 ^ w17135;
	assign w17210 = w46991 ^ w17137;
	assign w17213 = w46990 ^ w17137;
	assign w17212 = w17142 ^ w17137;
	assign w8733 = w8734 ^ w8735;
	assign w49532 = ~w8733;
	assign w46979 = w49532 ^ w944;
	assign w17001 = w46979 ^ w46977;
	assign w17018 = w46979 ^ w46978;
	assign w17003 = w46978 ^ w17001;
	assign w17078 = w17008 ^ w17003;
	assign w17079 = w46974 ^ w17003;
	assign w16554 = w46880 ^ w46877;
	assign w16546 = w16465 ^ w16554;
	assign w16545 = w46884 ^ w16546;
	assign w17076 = w46975 ^ w17003;
	assign w17084 = w46979 ^ w17088;
	assign w17071 = w17088 & w17084;
	assign w17924 = w17928 ^ w44125;
	assign w17923 = w17947 ^ w17924;
	assign w49699 = w17922 ^ w17923;
	assign w8829 = w49699 ^ w49704;
	assign w8774 = w8829 ^ w8815;
	assign w8557 = w8801 ^ w49699;
	assign w8877 = w8557 ^ w8558;
	assign w8750 = w8829 ^ w8819;
	assign w49637 = w49708 ^ w8750;
	assign w49621 = w49699 ^ w8775;
	assign w8762 = w8829 ^ w49712;
	assign w49629 = w8762 ^ w8763;
	assign w46874 = w49637 ^ w1877;
	assign w30224 = w46874 ^ w46872;
	assign w30221 = w46869 ^ w46874;
	assign w46890 = w49621 ^ w1861;
	assign w33303 = w46885 ^ w46890;
	assign w8772 = ~w8774;
	assign w46882 = w49629 ^ w1869;
	assign w16442 = w46881 ^ w46882;
	assign w16556 = w46882 ^ w46880;
	assign w16482 = w46883 ^ w46882;
	assign w16467 = w46882 ^ w16465;
	assign w16542 = w16472 ^ w16467;
	assign w16550 = w16554 ^ w16482;
	assign w16539 = w16546 & w16550;
	assign w16543 = w46878 ^ w16467;
	assign w16533 = w16554 & w16543;
	assign w16469 = w16533 ^ w16467;
	assign w16553 = w46877 ^ w46882;
	assign w16471 = w16539 ^ w16468;
	assign w16475 = w16471 ^ w16469;
	assign w16480 = w46877 ^ w16475;
	assign w17927 = w17966 ^ w17924;
	assign w18031 = w17926 ^ w17927;
	assign w45393 = ~w18031;
	assign w8768 = w18032 ^ w45393;
	assign w8766 = w8767 ^ w8768;
	assign w49625 = ~w8766;
	assign w49640 = w45393 ^ w8746;
	assign w8824 = w45393 ^ w45372;
	assign w8771 = w8855 ^ w8824;
	assign w8782 = w8824 ^ w8812;
	assign w49624 = w45380 ^ w8771;
	assign w46887 = w49624 ^ w1864;
	assign w33216 = w46887 ^ w46885;
	assign w46871 = w49640 ^ w1880;
	assign w30134 = w46871 ^ w46869;
	assign w30209 = w30134 ^ w30224;
	assign w30217 = w30134 ^ w30140;
	assign w30220 = w46871 ^ w30140;
	assign w30096 = w30136 ^ w30134;
	assign w30095 = w30136 ^ w46871;
	assign w30219 = w46876 ^ w30095;
	assign w30205 = w46876 & w30219;
	assign w30200 = w30224 & w30209;
	assign w49617 = w45774 ^ w8782;
	assign w46894 = w49617 ^ w1857;
	assign w16606 = w46900 ^ w46894;
	assign w16602 = w46896 ^ w46894;
	assign w16686 = w46895 ^ w16606;
	assign w16682 = w46899 ^ w16686;
	assign w16561 = w16602 ^ w46895;
	assign w16669 = w16686 & w16682;
	assign w46886 = w49625 ^ w1865;
	assign w33222 = w46892 ^ w46886;
	assign w33299 = w33216 ^ w33222;
	assign w33302 = w46887 ^ w33222;
	assign w8758 = w8824 ^ w49710;
	assign w49632 = w8758 ^ w8759;
	assign w46879 = w49632 ^ w1872;
	assign w16466 = w46879 ^ w46877;
	assign w16552 = w46879 ^ w16472;
	assign w16548 = w46883 ^ w16552;
	assign w16427 = w16468 ^ w46879;
	assign w16551 = w46884 ^ w16427;
	assign w16537 = w46884 & w16551;
	assign w16535 = w16552 & w16548;
	assign w16428 = w16468 ^ w16466;
	assign w16544 = w16465 ^ w16428;
	assign w16531 = w16553 & w16544;
	assign w16541 = w16466 ^ w16556;
	assign w16532 = w16556 & w16541;
	assign w16441 = w16532 ^ w16533;
	assign w16488 = w16441 ^ w16442;
	assign w16549 = w16466 ^ w16472;
	assign w16534 = w16549 & w16542;
	assign w44058 = w16531 ^ w16534;
	assign w16484 = w16532 ^ w44058;
	assign w16440 = w16535 ^ w16484;
	assign w16522 = w46883 ^ w16440;
	assign w16547 = w16482 ^ w16549;
	assign w16538 = w16547 & w16545;
	assign w16489 = w16532 ^ w16538;
	assign w16530 = w16489 ^ w16480;
	assign w44061 = w16531 ^ w16537;
	assign w16481 = w44061 ^ w16466;
	assign w16527 = w16489 ^ w16481;
	assign w16443 = w16475 ^ w44061;
	assign w16486 = w46879 ^ w16443;
	assign w16540 = w46879 ^ w16467;
	assign w16536 = w16555 & w16540;
	assign w16470 = w16536 ^ w16466;
	assign w16487 = w16488 ^ w16470;
	assign w16529 = w16535 ^ w16487;
	assign w16526 = w16530 & w16529;
	assign w16521 = w16526 ^ w16486;
	assign w16520 = w16521 & w16522;
	assign w16518 = w16526 ^ w16520;
	assign w16438 = w16520 ^ w16537;
	assign w16433 = w16438 ^ w16534;
	assign w16444 = w16470 ^ w44058;
	assign w16528 = w16444 ^ w16469;
	assign w16519 = w16520 ^ w16528;
	assign w16525 = w16526 ^ w16528;
	assign w16505 = w16519 & w46884;
	assign w16524 = w16527 & w16525;
	assign w16435 = w16524 ^ w16536;
	assign w16523 = w16524 ^ w16486;
	assign w16431 = w16435 ^ w16471;
	assign w16434 = w46877 ^ w16431;
	assign w16511 = w16433 ^ w16434;
	assign w16502 = w16523 & w16542;
	assign w16430 = w46879 ^ w16431;
	assign w16501 = w16511 & w16543;
	assign w16496 = w16519 & w16551;
	assign w16517 = w16528 & w16518;
	assign w16515 = w16517 ^ w16525;
	assign w16514 = w16523 & w16515;
	assign w16479 = w16514 ^ w16489;
	assign w16513 = w16479 ^ w16481;
	assign w16437 = w16514 ^ w16538;
	assign w16503 = w16513 & w16552;
	assign w16446 = w16502 ^ w16503;
	assign w16494 = w16513 & w16548;
	assign w16464 = w16502 ^ w16494;
	assign w16493 = w16523 & w16549;
	assign w16492 = w16511 & w16554;
	assign w44060 = w16517 ^ w16535;
	assign w16509 = w44060 ^ w16487;
	assign w16498 = w16509 & w16550;
	assign w16507 = w16509 & w16546;
	assign w16476 = w46883 ^ w44060;
	assign w44063 = w16505 ^ w16507;
	assign w16439 = w16520 ^ w16484;
	assign w16516 = w16476 ^ w16439;
	assign w16506 = w16516 & w16545;
	assign w16497 = w16516 & w16547;
	assign w16429 = w16476 ^ w16437;
	assign w16508 = w16429 ^ w16430;
	assign w16491 = w16508 & w16556;
	assign w16500 = w16508 & w16541;
	assign w16461 = w16500 ^ w16503;
	assign w16457 = w16500 ^ w16501;
	assign w16458 = ~w16461;
	assign w44059 = w16491 ^ w16492;
	assign w16473 = w16497 ^ w44059;
	assign w16474 = w16498 ^ w16473;
	assign w16478 = w16506 ^ w16474;
	assign w16483 = w16507 ^ w16478;
	assign w16558 = w16483 ^ w16457;
	assign w16447 = w16505 ^ w16478;
	assign w49856 = w16446 ^ w16447;
	assign w16460 = w16464 ^ w44059;
	assign w16436 = w16466 ^ w16429;
	assign w16512 = w16433 ^ w16436;
	assign w16499 = w16512 & w16544;
	assign w16490 = w16512 & w16553;
	assign w16456 = w16501 ^ w16490;
	assign w16452 = ~w16456;
	assign w16432 = w16524 ^ w16480;
	assign w16510 = w16479 ^ w16432;
	assign w16504 = w16510 & w16540;
	assign w16495 = w16510 & w16555;
	assign w16477 = w16495 ^ w16499;
	assign w16455 = ~w16477;
	assign w16462 = w16504 ^ w16495;
	assign w16454 = w16455 ^ w16493;
	assign w16450 = w16454 ^ w44063;
	assign w16453 = w16492 ^ w16450;
	assign w16449 = w16473 ^ w16450;
	assign w44062 = w16503 ^ w16504;
	assign w49857 = w44062 ^ w16483;
	assign w16485 = w16500 ^ w44062;
	assign w16451 = w16496 ^ w16485;
	assign w16445 = w16501 ^ w16485;
	assign w16448 = ~w16451;
	assign w49855 = w16448 ^ w16449;
	assign w49858 = w16474 ^ w16445;
	assign w9179 = w49848 ^ w49855;
	assign w9141 = w49853 ^ w49858;
	assign w8936 = ~w49855;
	assign w9114 = w45611 ^ w8936;
	assign w8935 = w49856 ^ w8936;
	assign w9075 = ~w9141;
	assign w9079 = w9075 ^ w45240;
	assign w9062 = ~w9179;
	assign w9073 = w9204 ^ w9062;
	assign w9060 = w9062 ^ w49844;
	assign w8927 = w49856 ^ w49849;
	assign w45348 = ~w16558;
	assign w9065 = w45348 ^ w12002;
	assign w16685 = w46900 ^ w16561;
	assign w16671 = w46900 & w16685;
	assign w9069 = w49857 ^ w49850;
	assign w16463 = w44063 ^ w16460;
	assign w16560 = w16462 ^ w16463;
	assign w45349 = ~w16560;
	assign w9180 = w45241 ^ w45349;
	assign w8933 = w45611 ^ w45349;
	assign w16459 = w16455 ^ w16460;
	assign w16559 = w16458 ^ w16459;
	assign w49854 = ~w16559;
	assign w9181 = w45240 ^ w49854;
	assign w8929 = w16559 ^ w45612;
	assign w16557 = w16452 ^ w16453;
	assign w45347 = ~w16557;
	assign w9067 = w45347 ^ w12001;
	assign w49614 = w8877 ^ w8809;
	assign w46897 = w49614 ^ w1854;
	assign w16599 = w46899 ^ w46897;
	assign w16601 = w46898 ^ w16599;
	assign w16676 = w16606 ^ w16601;
	assign w16677 = w46894 ^ w16601;
	assign w16674 = w46895 ^ w16601;
	assign w16576 = w46897 ^ w46898;
	assign w45933 = ~w8791;
	assign w8613 = w45933 ^ w45378;
	assign w49604 = w8612 ^ w8613;
	assign w46907 = w49604 ^ w888;
	assign w30350 = w46907 ^ w30354;
	assign w30284 = w46907 ^ w46906;
	assign w30349 = w30284 ^ w30351;
	assign w30357 = w46901 ^ w46907;
	assign w30337 = w30354 & w30350;
	assign w8608 = w45933 ^ w49692;
	assign w49606 = w8607 ^ w8608;
	assign w46905 = w49606 ^ w890;
	assign w30267 = w46907 ^ w46905;
	assign w30269 = w46906 ^ w30267;
	assign w30345 = w46902 ^ w30269;
	assign w30342 = w46903 ^ w30269;
	assign w30344 = w30274 ^ w30269;
	assign w30244 = w46905 ^ w46906;
	assign w30338 = w30357 & w30342;
	assign w30272 = w30338 ^ w30268;
	assign w30336 = w30351 & w30344;
	assign w8605 = w45933 ^ w49693;
	assign w49607 = w8604 ^ w8605;
	assign w46904 = w49607 ^ w891;
	assign w30270 = w46904 ^ w46902;
	assign w30356 = w46904 ^ w46901;
	assign w30352 = w30356 ^ w30284;
	assign w30348 = w30267 ^ w30356;
	assign w30347 = w46908 ^ w30348;
	assign w30358 = w46906 ^ w46904;
	assign w30343 = w30268 ^ w30358;
	assign w30230 = w30270 ^ w30268;
	assign w30346 = w30267 ^ w30230;
	assign w30229 = w30270 ^ w46903;
	assign w30353 = w46908 ^ w30229;
	assign w30341 = w30348 & w30352;
	assign w30273 = w30341 ^ w30270;
	assign w30340 = w30349 & w30347;
	assign w30339 = w46908 & w30353;
	assign w30335 = w30356 & w30345;
	assign w30271 = w30335 ^ w30269;
	assign w30277 = w30273 ^ w30271;
	assign w30282 = w46901 ^ w30277;
	assign w30334 = w30358 & w30343;
	assign w30291 = w30334 ^ w30340;
	assign w30332 = w30291 ^ w30282;
	assign w30243 = w30334 ^ w30335;
	assign w30290 = w30243 ^ w30244;
	assign w30289 = w30290 ^ w30272;
	assign w30331 = w30337 ^ w30289;
	assign w30333 = w30355 & w30346;
	assign w30328 = w30332 & w30331;
	assign w44637 = w30333 ^ w30339;
	assign w30245 = w30277 ^ w44637;
	assign w30288 = w46903 ^ w30245;
	assign w30323 = w30328 ^ w30288;
	assign w30283 = w44637 ^ w30268;
	assign w30329 = w30291 ^ w30283;
	assign w44638 = w30333 ^ w30336;
	assign w30286 = w30334 ^ w44638;
	assign w30242 = w30337 ^ w30286;
	assign w30324 = w46907 ^ w30242;
	assign w30322 = w30323 & w30324;
	assign w30241 = w30322 ^ w30286;
	assign w30320 = w30328 ^ w30322;
	assign w30240 = w30322 ^ w30339;
	assign w30235 = w30240 ^ w30336;
	assign w30246 = w30272 ^ w44638;
	assign w30330 = w30246 ^ w30271;
	assign w30321 = w30322 ^ w30330;
	assign w30327 = w30328 ^ w30330;
	assign w30326 = w30329 & w30327;
	assign w30325 = w30326 ^ w30288;
	assign w30237 = w30326 ^ w30338;
	assign w30233 = w30237 ^ w30273;
	assign w30236 = w46901 ^ w30233;
	assign w30313 = w30235 ^ w30236;
	assign w30234 = w30326 ^ w30282;
	assign w30232 = w46903 ^ w30233;
	assign w30319 = w30330 & w30320;
	assign w30317 = w30319 ^ w30327;
	assign w30316 = w30325 & w30317;
	assign w30281 = w30316 ^ w30291;
	assign w30315 = w30281 ^ w30283;
	assign w30239 = w30316 ^ w30340;
	assign w30312 = w30281 ^ w30234;
	assign w30307 = w30321 & w46908;
	assign w30306 = w30312 & w30342;
	assign w30305 = w30315 & w30354;
	assign w30304 = w30325 & w30344;
	assign w30248 = w30304 ^ w30305;
	assign w30303 = w30313 & w30345;
	assign w30298 = w30321 & w30353;
	assign w30297 = w30312 & w30357;
	assign w30264 = w30306 ^ w30297;
	assign w30296 = w30315 & w30350;
	assign w30266 = w30304 ^ w30296;
	assign w30295 = w30325 & w30351;
	assign w30294 = w30313 & w30356;
	assign w44640 = w30305 ^ w30306;
	assign w44642 = w30319 ^ w30337;
	assign w30311 = w44642 ^ w30289;
	assign w30309 = w30311 & w30348;
	assign w44641 = w30307 ^ w30309;
	assign w30300 = w30311 & w30352;
	assign w30278 = w46907 ^ w44642;
	assign w30318 = w30278 ^ w30241;
	assign w30231 = w30278 ^ w30239;
	assign w30238 = w30268 ^ w30231;
	assign w30314 = w30235 ^ w30238;
	assign w30310 = w30231 ^ w30232;
	assign w30308 = w30318 & w30347;
	assign w30302 = w30310 & w30343;
	assign w30287 = w30302 ^ w44640;
	assign w30263 = w30302 ^ w30305;
	assign w30260 = ~w30263;
	assign w30259 = w30302 ^ w30303;
	assign w30253 = w30298 ^ w30287;
	assign w30250 = ~w30253;
	assign w30247 = w30303 ^ w30287;
	assign w30301 = w30314 & w30346;
	assign w30279 = w30297 ^ w30301;
	assign w30257 = ~w30279;
	assign w30256 = w30257 ^ w30295;
	assign w30252 = w30256 ^ w44641;
	assign w30255 = w30294 ^ w30252;
	assign w30299 = w30318 & w30349;
	assign w30293 = w30310 & w30358;
	assign w30292 = w30314 & w30355;
	assign w30258 = w30303 ^ w30292;
	assign w30254 = ~w30258;
	assign w30359 = w30254 ^ w30255;
	assign w44639 = w30293 ^ w30294;
	assign w30275 = w30299 ^ w44639;
	assign w30251 = w30275 ^ w30252;
	assign w49896 = w30250 ^ w30251;
	assign w30276 = w30300 ^ w30275;
	assign w49899 = w30276 ^ w30247;
	assign w30280 = w30308 ^ w30276;
	assign w30249 = w30307 ^ w30280;
	assign w49897 = w30248 ^ w30249;
	assign w30285 = w30309 ^ w30280;
	assign w30360 = w30285 ^ w30259;
	assign w9135 = w49895 ^ w49899;
	assign w9175 = w49893 ^ w49897;
	assign w9185 = w49892 ^ w49896;
	assign w8998 = ~w9185;
	assign w49898 = w44640 ^ w30285;
	assign w9166 = w49894 ^ w49898;
	assign w30262 = w30266 ^ w44639;
	assign w30265 = w44641 ^ w30262;
	assign w30362 = w30264 ^ w30265;
	assign w30261 = w30257 ^ w30262;
	assign w30361 = w30260 ^ w30261;
	assign w45694 = ~w30359;
	assign w9160 = w45359 ^ w45694;
	assign w8995 = w9160 ^ w49898;
	assign w8993 = ~w8995;
	assign w45695 = ~w30360;
	assign w9149 = w45360 ^ w45695;
	assign w8985 = w9135 ^ w45695;
	assign w8988 = w9149 ^ w45694;
	assign w45696 = ~w30361;
	assign w9189 = w45361 ^ w45696;
	assign w8996 = w8998 ^ w45696;
	assign w45697 = ~w30362;
	assign w9197 = w45354 ^ w45697;
	assign w45934 = ~w8790;
	assign w8593 = w45934 ^ w49700;
	assign w8862 = w8593 ^ w8594;
	assign w49623 = w8862 ^ w8806;
	assign w46888 = w49623 ^ w1863;
	assign w33218 = w46888 ^ w46886;
	assign w33304 = w46888 ^ w46885;
	assign w33306 = w46890 ^ w46888;
	assign w33291 = w33216 ^ w33306;
	assign w33178 = w33218 ^ w33216;
	assign w33177 = w33218 ^ w46887;
	assign w33301 = w46892 ^ w33177;
	assign w33287 = w46892 & w33301;
	assign w33282 = w33306 & w33291;
	assign w8778 = w45934 ^ w45386;
	assign w8776 = w8777 ^ w8778;
	assign w49620 = ~w8776;
	assign w46891 = w49620 ^ w1860;
	assign w33298 = w46891 ^ w33302;
	assign w33232 = w46891 ^ w46890;
	assign w33297 = w33232 ^ w33299;
	assign w33300 = w33304 ^ w33232;
	assign w33305 = w46885 ^ w46891;
	assign w33285 = w33302 & w33298;
	assign w8773 = w45934 ^ w49709;
	assign w49622 = w8772 ^ w8773;
	assign w46889 = w49622 ^ w1862;
	assign w33215 = w46891 ^ w46889;
	assign w33217 = w46890 ^ w33215;
	assign w33293 = w46886 ^ w33217;
	assign w33290 = w46887 ^ w33217;
	assign w33292 = w33222 ^ w33217;
	assign w33296 = w33215 ^ w33304;
	assign w33295 = w46892 ^ w33296;
	assign w33192 = w46889 ^ w46890;
	assign w33294 = w33215 ^ w33178;
	assign w33289 = w33296 & w33300;
	assign w33221 = w33289 ^ w33218;
	assign w33288 = w33297 & w33295;
	assign w33239 = w33282 ^ w33288;
	assign w33286 = w33305 & w33290;
	assign w33220 = w33286 ^ w33216;
	assign w33284 = w33299 & w33292;
	assign w33283 = w33304 & w33293;
	assign w33219 = w33283 ^ w33217;
	assign w33225 = w33221 ^ w33219;
	assign w33230 = w46885 ^ w33225;
	assign w33280 = w33239 ^ w33230;
	assign w33191 = w33282 ^ w33283;
	assign w33238 = w33191 ^ w33192;
	assign w33237 = w33238 ^ w33220;
	assign w33279 = w33285 ^ w33237;
	assign w33281 = w33303 & w33294;
	assign w33276 = w33280 & w33279;
	assign w44760 = w33281 ^ w33287;
	assign w33193 = w33225 ^ w44760;
	assign w33236 = w46887 ^ w33193;
	assign w33271 = w33276 ^ w33236;
	assign w33231 = w44760 ^ w33216;
	assign w33277 = w33239 ^ w33231;
	assign w44761 = w33281 ^ w33284;
	assign w33234 = w33282 ^ w44761;
	assign w33190 = w33285 ^ w33234;
	assign w33272 = w46891 ^ w33190;
	assign w33270 = w33271 & w33272;
	assign w33189 = w33270 ^ w33234;
	assign w33268 = w33276 ^ w33270;
	assign w33188 = w33270 ^ w33287;
	assign w33183 = w33188 ^ w33284;
	assign w33194 = w33220 ^ w44761;
	assign w33278 = w33194 ^ w33219;
	assign w33269 = w33270 ^ w33278;
	assign w33275 = w33276 ^ w33278;
	assign w33274 = w33277 & w33275;
	assign w33273 = w33274 ^ w33236;
	assign w33185 = w33274 ^ w33286;
	assign w33181 = w33185 ^ w33221;
	assign w33184 = w46885 ^ w33181;
	assign w33261 = w33183 ^ w33184;
	assign w33182 = w33274 ^ w33230;
	assign w33180 = w46887 ^ w33181;
	assign w33267 = w33278 & w33268;
	assign w33265 = w33267 ^ w33275;
	assign w33264 = w33273 & w33265;
	assign w33229 = w33264 ^ w33239;
	assign w33263 = w33229 ^ w33231;
	assign w33187 = w33264 ^ w33288;
	assign w33260 = w33229 ^ w33182;
	assign w33255 = w33269 & w46892;
	assign w33254 = w33260 & w33290;
	assign w33253 = w33263 & w33302;
	assign w33252 = w33273 & w33292;
	assign w33196 = w33252 ^ w33253;
	assign w33251 = w33261 & w33293;
	assign w33246 = w33269 & w33301;
	assign w33245 = w33260 & w33305;
	assign w33212 = w33254 ^ w33245;
	assign w33244 = w33263 & w33298;
	assign w33214 = w33252 ^ w33244;
	assign w33243 = w33273 & w33299;
	assign w33242 = w33261 & w33304;
	assign w44763 = w33253 ^ w33254;
	assign w44765 = w33267 ^ w33285;
	assign w33259 = w44765 ^ w33237;
	assign w33257 = w33259 & w33296;
	assign w44764 = w33255 ^ w33257;
	assign w33248 = w33259 & w33300;
	assign w33226 = w46891 ^ w44765;
	assign w33266 = w33226 ^ w33189;
	assign w33179 = w33226 ^ w33187;
	assign w33186 = w33216 ^ w33179;
	assign w33262 = w33183 ^ w33186;
	assign w33258 = w33179 ^ w33180;
	assign w33256 = w33266 & w33295;
	assign w33250 = w33258 & w33291;
	assign w33235 = w33250 ^ w44763;
	assign w33211 = w33250 ^ w33253;
	assign w33208 = ~w33211;
	assign w33207 = w33250 ^ w33251;
	assign w33201 = w33246 ^ w33235;
	assign w33198 = ~w33201;
	assign w33195 = w33251 ^ w33235;
	assign w33249 = w33262 & w33294;
	assign w33227 = w33245 ^ w33249;
	assign w33205 = ~w33227;
	assign w33204 = w33205 ^ w33243;
	assign w33200 = w33204 ^ w44764;
	assign w33203 = w33242 ^ w33200;
	assign w33247 = w33266 & w33297;
	assign w33241 = w33258 & w33306;
	assign w33240 = w33262 & w33303;
	assign w33206 = w33251 ^ w33240;
	assign w33202 = ~w33206;
	assign w33307 = w33202 ^ w33203;
	assign w44762 = w33241 ^ w33242;
	assign w33223 = w33247 ^ w44762;
	assign w33199 = w33223 ^ w33200;
	assign w49869 = w33198 ^ w33199;
	assign w33224 = w33248 ^ w33223;
	assign w49872 = w33224 ^ w33195;
	assign w33228 = w33256 ^ w33224;
	assign w33197 = w33255 ^ w33228;
	assign w49870 = w33196 ^ w33197;
	assign w33233 = w33257 ^ w33228;
	assign w33308 = w33233 ^ w33207;
	assign w9137 = w49867 ^ w49872;
	assign w9169 = w49865 ^ w49870;
	assign w9172 = w49864 ^ w49869;
	assign w9000 = w9137 ^ w45523;
	assign w9025 = ~w9172;
	assign w9033 = ~w9169;
	assign w9023 = w9025 ^ w49877;
	assign w8896 = ~w49870;
	assign w8895 = w8896 ^ w49864;
	assign w9224 = w8894 ^ w8895;
	assign w49871 = w44763 ^ w33233;
	assign w9165 = w49866 ^ w49871;
	assign w9007 = ~w9165;
	assign w33210 = w33214 ^ w44762;
	assign w33213 = w44764 ^ w33210;
	assign w33310 = w33212 ^ w33213;
	assign w33209 = w33205 ^ w33210;
	assign w33309 = w33208 ^ w33209;
	assign w49868 = ~w33309;
	assign w9176 = w45357 ^ w49868;
	assign w8892 = w33309 ^ w45350;
	assign w9225 = w8891 ^ w8892;
	assign w9051 = w49869 ^ w45357;
	assign w8898 = w49871 ^ w49865;
	assign w9223 = w8897 ^ w8898;
	assign w45770 = ~w33307;
	assign w9161 = w45355 ^ w45770;
	assign w9049 = w45770 ^ w49866;
	assign w9029 = w9161 ^ w9155;
	assign w9022 = w9161 ^ w45522;
	assign w9020 = ~w9022;
	assign w45771 = ~w33308;
	assign w9019 = w45771 ^ w45770;
	assign w45772 = ~w33310;
	assign w9177 = w45350 ^ w45772;
	assign w45935 = ~w8789;
	assign w8749 = w45935 ^ w49700;
	assign w8747 = w8748 ^ w8749;
	assign w49638 = ~w8747;
	assign w8752 = w45935 ^ w45374;
	assign w49636 = w8751 ^ w8752;
	assign w46873 = w49638 ^ w1878;
	assign w30110 = w46873 ^ w46874;
	assign w8780 = w45935 ^ w45373;
	assign w49618 = w8780 ^ w8781;
	assign w46893 = w49618 ^ w1858;
	assign w16600 = w46895 ^ w46893;
	assign w16675 = w16600 ^ w16690;
	assign w16683 = w16600 ^ w16606;
	assign w16681 = w16616 ^ w16683;
	assign w16562 = w16602 ^ w16600;
	assign w16689 = w46893 ^ w46899;
	assign w16670 = w16689 & w16674;
	assign w16604 = w16670 ^ w16600;
	assign w16687 = w46893 ^ w46898;
	assign w16666 = w16690 & w16675;
	assign w46875 = w49636 ^ w1876;
	assign w30133 = w46875 ^ w46873;
	assign w30135 = w46874 ^ w30133;
	assign w30211 = w46870 ^ w30135;
	assign w30208 = w46871 ^ w30135;
	assign w30210 = w30140 ^ w30135;
	assign w30216 = w46875 ^ w30220;
	assign w30214 = w30133 ^ w30222;
	assign w30213 = w46876 ^ w30214;
	assign w30150 = w46875 ^ w46874;
	assign w30215 = w30150 ^ w30217;
	assign w30218 = w30222 ^ w30150;
	assign w30212 = w30133 ^ w30096;
	assign w30223 = w46869 ^ w46875;
	assign w30207 = w30214 & w30218;
	assign w30139 = w30207 ^ w30136;
	assign w30206 = w30215 & w30213;
	assign w30157 = w30200 ^ w30206;
	assign w30204 = w30223 & w30208;
	assign w30138 = w30204 ^ w30134;
	assign w30203 = w30220 & w30216;
	assign w30202 = w30217 & w30210;
	assign w30201 = w30222 & w30211;
	assign w30137 = w30201 ^ w30135;
	assign w30143 = w30139 ^ w30137;
	assign w30148 = w46869 ^ w30143;
	assign w30198 = w30157 ^ w30148;
	assign w30109 = w30200 ^ w30201;
	assign w30156 = w30109 ^ w30110;
	assign w30155 = w30156 ^ w30138;
	assign w30197 = w30203 ^ w30155;
	assign w30199 = w30221 & w30212;
	assign w30194 = w30198 & w30197;
	assign w16678 = w16599 ^ w16562;
	assign w16665 = w16687 & w16678;
	assign w44064 = w16665 ^ w16671;
	assign w16615 = w44064 ^ w16600;
	assign w16668 = w16683 & w16676;
	assign w44065 = w16665 ^ w16668;
	assign w16618 = w16666 ^ w44065;
	assign w16574 = w16669 ^ w16618;
	assign w16656 = w46899 ^ w16574;
	assign w44632 = w30199 ^ w30205;
	assign w30149 = w44632 ^ w30134;
	assign w30195 = w30157 ^ w30149;
	assign w30111 = w30143 ^ w44632;
	assign w30154 = w46871 ^ w30111;
	assign w30189 = w30194 ^ w30154;
	assign w44633 = w30199 ^ w30202;
	assign w30152 = w30200 ^ w44633;
	assign w30108 = w30203 ^ w30152;
	assign w30190 = w46875 ^ w30108;
	assign w30188 = w30189 & w30190;
	assign w30107 = w30188 ^ w30152;
	assign w30106 = w30188 ^ w30205;
	assign w30101 = w30106 ^ w30202;
	assign w30186 = w30194 ^ w30188;
	assign w30112 = w30138 ^ w44633;
	assign w30196 = w30112 ^ w30137;
	assign w30187 = w30188 ^ w30196;
	assign w30193 = w30194 ^ w30196;
	assign w30192 = w30195 & w30193;
	assign w30191 = w30192 ^ w30154;
	assign w30103 = w30192 ^ w30204;
	assign w30099 = w30103 ^ w30139;
	assign w30102 = w46869 ^ w30099;
	assign w30179 = w30101 ^ w30102;
	assign w30100 = w30192 ^ w30148;
	assign w30098 = w46871 ^ w30099;
	assign w30185 = w30196 & w30186;
	assign w30183 = w30185 ^ w30193;
	assign w30182 = w30191 & w30183;
	assign w30147 = w30182 ^ w30157;
	assign w30181 = w30147 ^ w30149;
	assign w30105 = w30182 ^ w30206;
	assign w30178 = w30147 ^ w30100;
	assign w30173 = w30187 & w46876;
	assign w30172 = w30178 & w30208;
	assign w30171 = w30181 & w30220;
	assign w30170 = w30191 & w30210;
	assign w30114 = w30170 ^ w30171;
	assign w30169 = w30179 & w30211;
	assign w30164 = w30187 & w30219;
	assign w30163 = w30178 & w30223;
	assign w30130 = w30172 ^ w30163;
	assign w30162 = w30181 & w30216;
	assign w30132 = w30170 ^ w30162;
	assign w30161 = w30191 & w30217;
	assign w30160 = w30179 & w30222;
	assign w44634 = w30171 ^ w30172;
	assign w44636 = w30185 ^ w30203;
	assign w30144 = w46875 ^ w44636;
	assign w30184 = w30144 ^ w30107;
	assign w30165 = w30184 & w30215;
	assign w30174 = w30184 & w30213;
	assign w30097 = w30144 ^ w30105;
	assign w30104 = w30134 ^ w30097;
	assign w30180 = w30101 ^ w30104;
	assign w30167 = w30180 & w30212;
	assign w30145 = w30163 ^ w30167;
	assign w30123 = ~w30145;
	assign w30122 = w30123 ^ w30161;
	assign w30176 = w30097 ^ w30098;
	assign w30159 = w30176 & w30224;
	assign w30158 = w30180 & w30221;
	assign w30124 = w30169 ^ w30158;
	assign w30120 = ~w30124;
	assign w43583 = w30159 ^ w30160;
	assign w30128 = w30132 ^ w43583;
	assign w30127 = w30123 ^ w30128;
	assign w30141 = w30165 ^ w43583;
	assign w30168 = w30176 & w30209;
	assign w30125 = w30168 ^ w30169;
	assign w30153 = w30168 ^ w44634;
	assign w30119 = w30164 ^ w30153;
	assign w30116 = ~w30119;
	assign w30113 = w30169 ^ w30153;
	assign w30129 = w30168 ^ w30171;
	assign w30126 = ~w30129;
	assign w30227 = w30126 ^ w30127;
	assign w30177 = w44636 ^ w30155;
	assign w30175 = w30177 & w30214;
	assign w30166 = w30177 & w30218;
	assign w30142 = w30166 ^ w30141;
	assign w30146 = w30174 ^ w30142;
	assign w30151 = w30175 ^ w30146;
	assign w49915 = w44634 ^ w30151;
	assign w30226 = w30151 ^ w30125;
	assign w30115 = w30173 ^ w30146;
	assign w49914 = w30114 ^ w30115;
	assign w49916 = w30142 ^ w30113;
	assign w9150 = w49911 ^ w49915;
	assign w9133 = w49912 ^ w49916;
	assign w9229 = ~w9133;
	assign w9096 = w9229 ^ w45607;
	assign w44635 = w30173 ^ w30175;
	assign w30131 = w44635 ^ w30128;
	assign w30228 = w30130 ^ w30131;
	assign w30118 = w30122 ^ w44635;
	assign w30121 = w30160 ^ w30118;
	assign w30225 = w30120 ^ w30121;
	assign w30117 = w30141 ^ w30118;
	assign w49913 = w30116 ^ w30117;
	assign w9151 = w49909 ^ w49913;
	assign w8902 = w49914 ^ w49913;
	assign w16688 = w46896 ^ w46893;
	assign w16684 = w16688 ^ w16616;
	assign w16667 = w16688 & w16677;
	assign w16603 = w16667 ^ w16601;
	assign w16575 = w16666 ^ w16667;
	assign w16622 = w16575 ^ w16576;
	assign w16621 = w16622 ^ w16604;
	assign w16663 = w16669 ^ w16621;
	assign w16680 = w16599 ^ w16688;
	assign w16679 = w46900 ^ w16680;
	assign w16672 = w16681 & w16679;
	assign w16623 = w16666 ^ w16672;
	assign w16661 = w16623 ^ w16615;
	assign w16673 = w16680 & w16684;
	assign w16605 = w16673 ^ w16602;
	assign w16609 = w16605 ^ w16603;
	assign w16614 = w46893 ^ w16609;
	assign w16664 = w16623 ^ w16614;
	assign w16577 = w16609 ^ w44064;
	assign w16620 = w46895 ^ w16577;
	assign w16660 = w16664 & w16663;
	assign w16655 = w16660 ^ w16620;
	assign w16654 = w16655 & w16656;
	assign w16652 = w16660 ^ w16654;
	assign w16573 = w16654 ^ w16618;
	assign w16572 = w16654 ^ w16671;
	assign w16567 = w16572 ^ w16668;
	assign w16578 = w16604 ^ w44065;
	assign w16662 = w16578 ^ w16603;
	assign w16653 = w16654 ^ w16662;
	assign w16651 = w16662 & w16652;
	assign w16630 = w16653 & w16685;
	assign w16639 = w16653 & w46900;
	assign w16659 = w16660 ^ w16662;
	assign w16649 = w16651 ^ w16659;
	assign w16658 = w16661 & w16659;
	assign w16657 = w16658 ^ w16620;
	assign w16648 = w16657 & w16649;
	assign w16613 = w16648 ^ w16623;
	assign w16647 = w16613 ^ w16615;
	assign w16627 = w16657 & w16683;
	assign w16637 = w16647 & w16686;
	assign w16628 = w16647 & w16682;
	assign w16636 = w16657 & w16676;
	assign w16580 = w16636 ^ w16637;
	assign w16598 = w16636 ^ w16628;
	assign w16566 = w16658 ^ w16614;
	assign w16644 = w16613 ^ w16566;
	assign w16629 = w16644 & w16689;
	assign w16638 = w16644 & w16674;
	assign w16596 = w16638 ^ w16629;
	assign w44067 = w16637 ^ w16638;
	assign w44069 = w16651 ^ w16669;
	assign w16643 = w44069 ^ w16621;
	assign w16632 = w16643 & w16684;
	assign w16641 = w16643 & w16680;
	assign w44068 = w16639 ^ w16641;
	assign w16610 = w46899 ^ w44069;
	assign w16650 = w16610 ^ w16573;
	assign w16640 = w16650 & w16679;
	assign w16631 = w16650 & w16681;
	assign w16569 = w16658 ^ w16670;
	assign w16565 = w16569 ^ w16605;
	assign w16564 = w46895 ^ w16565;
	assign w8940 = w9133 ^ w49914;
	assign w9205 = w8940 ^ w8941;
	assign w45690 = ~w30225;
	assign w45691 = ~w30226;
	assign w9156 = w45606 ^ w45691;
	assign w9124 = w9229 ^ w45691;
	assign w45692 = ~w30227;
	assign w9163 = w45607 ^ w45692;
	assign w45693 = ~w30228;
	assign w9183 = w45608 ^ w45693;
	assign w16568 = w46893 ^ w16565;
	assign w16645 = w16567 ^ w16568;
	assign w16626 = w16645 & w16688;
	assign w16635 = w16645 & w16677;
	assign w16571 = w16648 ^ w16672;
	assign w16563 = w16610 ^ w16571;
	assign w16642 = w16563 ^ w16564;
	assign w16625 = w16642 & w16690;
	assign w16634 = w16642 & w16675;
	assign w16619 = w16634 ^ w44067;
	assign w16585 = w16630 ^ w16619;
	assign w16591 = w16634 ^ w16635;
	assign w16582 = ~w16585;
	assign w44066 = w16625 ^ w16626;
	assign w16607 = w16631 ^ w44066;
	assign w16608 = w16632 ^ w16607;
	assign w16612 = w16640 ^ w16608;
	assign w16617 = w16641 ^ w16612;
	assign w49883 = w44067 ^ w16617;
	assign w16581 = w16639 ^ w16612;
	assign w49882 = w16580 ^ w16581;
	assign w16594 = w16598 ^ w44066;
	assign w16579 = w16635 ^ w16619;
	assign w49884 = w16608 ^ w16579;
	assign w9143 = w49884 ^ w49899;
	assign w8999 = w9197 ^ w9143;
	assign w8912 = ~w9143;
	assign w8910 = w8912 ^ w45697;
	assign w8916 = w9143 ^ w49897;
	assign w8913 = w8912 ^ w49896;
	assign w16570 = w16600 ^ w16563;
	assign w16646 = w16567 ^ w16570;
	assign w16633 = w16646 & w16678;
	assign w16611 = w16629 ^ w16633;
	assign w16624 = w16646 & w16687;
	assign w16590 = w16635 ^ w16624;
	assign w16597 = w44068 ^ w16594;
	assign w16694 = w16596 ^ w16597;
	assign w45346 = ~w16694;
	assign w16595 = w16634 ^ w16637;
	assign w16592 = ~w16595;
	assign w16589 = ~w16611;
	assign w16593 = w16589 ^ w16594;
	assign w16693 = w16592 ^ w16593;
	assign w45353 = ~w16693;
	assign w16692 = w16617 ^ w16591;
	assign w45352 = ~w16692;
	assign w16586 = ~w16590;
	assign w16588 = w16589 ^ w16627;
	assign w16584 = w16588 ^ w44068;
	assign w16587 = w16626 ^ w16584;
	assign w16691 = w16586 ^ w16587;
	assign w16583 = w16607 ^ w16584;
	assign w49881 = w16582 ^ w16583;
	assign w45351 = ~w16691;
	assign w45936 = ~w8796;
	assign w8584 = w45936 ^ w45248;
	assign w8866 = w8584 ^ w8585;
	assign w8720 = w45936 ^ w49662;
	assign w49538 = w8720 ^ w8721;
	assign w46973 = w49538 ^ w950;
	assign w17090 = w46976 ^ w46973;
	assign w17086 = w17090 ^ w17018;
	assign w17069 = w17090 & w17079;
	assign w8741 = w45936 ^ w49645;
	assign w49527 = w8740 ^ w8741;
	assign w17002 = w46975 ^ w46973;
	assign w17077 = w17002 ^ w17092;
	assign w17068 = w17092 & w17077;
	assign w16964 = w17004 ^ w17002;
	assign w17080 = w17001 ^ w16964;
	assign w16977 = w17068 ^ w17069;
	assign w17085 = w17002 ^ w17008;
	assign w17070 = w17085 & w17078;
	assign w46984 = w49527 ^ w939;
	assign w33352 = w46984 ^ w46982;
	assign w33438 = w46984 ^ w46981;
	assign w33440 = w46986 ^ w46984;
	assign w33425 = w33350 ^ w33440;
	assign w33312 = w33352 ^ w33350;
	assign w33311 = w33352 ^ w46983;
	assign w33435 = w46988 ^ w33311;
	assign w33421 = w46988 & w33435;
	assign w33416 = w33440 & w33425;
	assign w17083 = w17018 ^ w17085;
	assign w17089 = w46973 ^ w46978;
	assign w17067 = w17089 & w17080;
	assign w17082 = w17001 ^ w17090;
	assign w17081 = w46980 ^ w17082;
	assign w17074 = w17083 & w17081;
	assign w17025 = w17068 ^ w17074;
	assign w17075 = w17082 & w17086;
	assign w17007 = w17075 ^ w17004;
	assign w44081 = w17067 ^ w17070;
	assign w17020 = w17068 ^ w44081;
	assign w16976 = w17071 ^ w17020;
	assign w17058 = w46979 ^ w16976;
	assign w44084 = w17067 ^ w17073;
	assign w17017 = w44084 ^ w17002;
	assign w17063 = w17025 ^ w17017;
	assign w49524 = w8866 ^ w8858;
	assign w46987 = w49524 ^ w936;
	assign w33349 = w46987 ^ w46985;
	assign w33351 = w46986 ^ w33349;
	assign w33427 = w46982 ^ w33351;
	assign w33424 = w46983 ^ w33351;
	assign w33426 = w33356 ^ w33351;
	assign w33432 = w46987 ^ w33436;
	assign w33430 = w33349 ^ w33438;
	assign w33429 = w46988 ^ w33430;
	assign w33366 = w46987 ^ w46986;
	assign w33431 = w33366 ^ w33433;
	assign w33434 = w33438 ^ w33366;
	assign w33428 = w33349 ^ w33312;
	assign w33439 = w46981 ^ w46987;
	assign w33423 = w33430 & w33434;
	assign w33355 = w33423 ^ w33352;
	assign w33422 = w33431 & w33429;
	assign w33373 = w33416 ^ w33422;
	assign w33420 = w33439 & w33424;
	assign w33354 = w33420 ^ w33350;
	assign w33419 = w33436 & w33432;
	assign w33418 = w33433 & w33426;
	assign w33417 = w33438 & w33427;
	assign w33353 = w33417 ^ w33351;
	assign w33359 = w33355 ^ w33353;
	assign w33364 = w46981 ^ w33359;
	assign w33414 = w33373 ^ w33364;
	assign w33325 = w33416 ^ w33417;
	assign w33372 = w33325 ^ w33326;
	assign w33371 = w33372 ^ w33354;
	assign w33413 = w33419 ^ w33371;
	assign w33415 = w33437 & w33428;
	assign w33410 = w33414 & w33413;
	assign w44766 = w33415 ^ w33421;
	assign w33365 = w44766 ^ w33350;
	assign w33411 = w33373 ^ w33365;
	assign w33327 = w33359 ^ w44766;
	assign w33370 = w46983 ^ w33327;
	assign w33405 = w33410 ^ w33370;
	assign w44767 = w33415 ^ w33418;
	assign w33368 = w33416 ^ w44767;
	assign w33324 = w33419 ^ w33368;
	assign w33406 = w46987 ^ w33324;
	assign w33404 = w33405 & w33406;
	assign w33323 = w33404 ^ w33368;
	assign w33322 = w33404 ^ w33421;
	assign w33317 = w33322 ^ w33418;
	assign w33402 = w33410 ^ w33404;
	assign w33328 = w33354 ^ w44767;
	assign w33412 = w33328 ^ w33353;
	assign w33403 = w33404 ^ w33412;
	assign w33409 = w33410 ^ w33412;
	assign w33408 = w33411 & w33409;
	assign w33407 = w33408 ^ w33370;
	assign w33319 = w33408 ^ w33420;
	assign w33315 = w33319 ^ w33355;
	assign w33318 = w46981 ^ w33315;
	assign w33395 = w33317 ^ w33318;
	assign w33316 = w33408 ^ w33364;
	assign w33314 = w46983 ^ w33315;
	assign w33401 = w33412 & w33402;
	assign w33399 = w33401 ^ w33409;
	assign w33398 = w33407 & w33399;
	assign w33363 = w33398 ^ w33373;
	assign w33397 = w33363 ^ w33365;
	assign w33321 = w33398 ^ w33422;
	assign w33394 = w33363 ^ w33316;
	assign w33389 = w33403 & w46988;
	assign w33388 = w33394 & w33424;
	assign w33387 = w33397 & w33436;
	assign w33386 = w33407 & w33426;
	assign w33330 = w33386 ^ w33387;
	assign w33385 = w33395 & w33427;
	assign w33380 = w33403 & w33435;
	assign w33379 = w33394 & w33439;
	assign w33346 = w33388 ^ w33379;
	assign w33378 = w33397 & w33432;
	assign w33348 = w33386 ^ w33378;
	assign w33377 = w33407 & w33433;
	assign w33376 = w33395 & w33438;
	assign w44768 = w33387 ^ w33388;
	assign w44770 = w33401 ^ w33419;
	assign w33360 = w46987 ^ w44770;
	assign w33400 = w33360 ^ w33323;
	assign w33381 = w33400 & w33431;
	assign w33390 = w33400 & w33429;
	assign w33313 = w33360 ^ w33321;
	assign w33320 = w33350 ^ w33313;
	assign w33396 = w33317 ^ w33320;
	assign w33383 = w33396 & w33428;
	assign w33361 = w33379 ^ w33383;
	assign w33339 = ~w33361;
	assign w33338 = w33339 ^ w33377;
	assign w33392 = w33313 ^ w33314;
	assign w33375 = w33392 & w33440;
	assign w33374 = w33396 & w33437;
	assign w33340 = w33385 ^ w33374;
	assign w33336 = ~w33340;
	assign w43593 = w33375 ^ w33376;
	assign w33344 = w33348 ^ w43593;
	assign w33343 = w33339 ^ w33344;
	assign w33357 = w33381 ^ w43593;
	assign w33384 = w33392 & w33425;
	assign w33341 = w33384 ^ w33385;
	assign w33369 = w33384 ^ w44768;
	assign w33335 = w33380 ^ w33369;
	assign w33332 = ~w33335;
	assign w33329 = w33385 ^ w33369;
	assign w33345 = w33384 ^ w33387;
	assign w33342 = ~w33345;
	assign w33443 = w33342 ^ w33343;
	assign w8911 = w33443 ^ w45346;
	assign w9217 = w8910 ^ w8911;
	assign w49781 = w9217 ^ w9189;
	assign w49885 = ~w33443;
	assign w46803 = w49781 ^ w991;
	assign w9200 = w45353 ^ w49885;
	assign w8958 = w9200 ^ w9197;
	assign w8956 = ~w8958;
	assign w8968 = w45361 ^ w33443;
	assign w8980 = w9200 ^ w9185;
	assign w49790 = w49881 ^ w8980;
	assign w46794 = w49790 ^ w1000;
	assign w33393 = w44770 ^ w33371;
	assign w33391 = w33393 & w33430;
	assign w33382 = w33393 & w33434;
	assign w33358 = w33382 ^ w33357;
	assign w33362 = w33390 ^ w33358;
	assign w33367 = w33391 ^ w33362;
	assign w49888 = w44768 ^ w33367;
	assign w33442 = w33367 ^ w33341;
	assign w33331 = w33389 ^ w33362;
	assign w49887 = w33330 ^ w33331;
	assign w49891 = w33358 ^ w33329;
	assign w49890 = ~w33442;
	assign w9142 = w49891 ^ w49895;
	assign w9164 = w45352 ^ w49890;
	assign w8973 = w9164 ^ w9135;
	assign w49795 = w49884 ^ w8973;
	assign w46789 = w49795 ^ w1005;
	assign w33169 = w46789 ^ w46794;
	assign w9178 = w49883 ^ w49888;
	assign w8950 = ~w9178;
	assign w8948 = w8950 ^ w9175;
	assign w9186 = w49882 ^ w49887;
	assign w8953 = ~w9186;
	assign w8951 = w8953 ^ w9185;
	assign w8961 = w45360 ^ w33442;
	assign w8976 = w8953 ^ w9166;
	assign w8986 = w49891 ^ w45352;
	assign w8964 = w9164 ^ w45695;
	assign w8962 = ~w8964;
	assign w8989 = w33442 ^ w45351;
	assign w8987 = w8988 ^ w8989;
	assign w49786 = ~w8987;
	assign w46798 = w49786 ^ w996;
	assign w49787 = w8985 ^ w8986;
	assign w46797 = w49787 ^ w997;
	assign w16153 = w46797 ^ w46803;
	assign w8975 = w9178 ^ w9160;
	assign w49793 = w45351 ^ w8975;
	assign w46791 = w49793 ^ w1003;
	assign w33082 = w46791 ^ w46789;
	assign w8917 = w49888 ^ w49882;
	assign w9215 = w8916 ^ w8917;
	assign w49784 = w9215 ^ w9166;
	assign w46800 = w49784 ^ w994;
	assign w16066 = w46800 ^ w46798;
	assign w16152 = w46800 ^ w46797;
	assign w8915 = ~w49887;
	assign w8914 = w8915 ^ w49881;
	assign w9216 = w8913 ^ w8914;
	assign w49783 = w9216 ^ w9175;
	assign w46801 = w49783 ^ w993;
	assign w16063 = w46803 ^ w46801;
	assign w16144 = w16063 ^ w16152;
	assign w8923 = ~w9142;
	assign w8924 = w8923 ^ w49898;
	assign w8920 = w8923 ^ w49897;
	assign w8918 = w9142 ^ w45696;
	assign w8925 = w49893 ^ w8915;
	assign w9212 = w8924 ^ w8925;
	assign w49800 = w9212 ^ w9178;
	assign w46784 = w49800 ^ w1010;
	assign w44769 = w33389 ^ w33391;
	assign w33347 = w44769 ^ w33344;
	assign w33444 = w33346 ^ w33347;
	assign w33334 = w33338 ^ w44769;
	assign w33337 = w33376 ^ w33334;
	assign w33441 = w33336 ^ w33337;
	assign w33333 = w33357 ^ w33334;
	assign w49886 = w33332 ^ w33333;
	assign w49889 = ~w33441;
	assign w9171 = w45351 ^ w49889;
	assign w8963 = w45359 ^ w33441;
	assign w49802 = w8962 ^ w8963;
	assign w46782 = w49802 ^ w1012;
	assign w8974 = w9171 ^ w9149;
	assign w8965 = w9171 ^ w45694;
	assign w8922 = ~w49886;
	assign w8997 = w8922 ^ w45353;
	assign w49782 = w8996 ^ w8997;
	assign w46802 = w49782 ^ w992;
	assign w16065 = w46802 ^ w16063;
	assign w16151 = w46797 ^ w46802;
	assign w16141 = w46798 ^ w16065;
	assign w16080 = w46803 ^ w46802;
	assign w16131 = w16152 & w16141;
	assign w16067 = w16131 ^ w16065;
	assign w16148 = w16152 ^ w16080;
	assign w16137 = w16144 & w16148;
	assign w16069 = w16137 ^ w16066;
	assign w16073 = w16069 ^ w16067;
	assign w16078 = w46797 ^ w16073;
	assign w16154 = w46802 ^ w46800;
	assign w9193 = w49881 ^ w49886;
	assign w8954 = w9193 ^ w9189;
	assign w49806 = w49892 ^ w8954;
	assign w46778 = w49806 ^ w1016;
	assign w8994 = w33441 ^ w49883;
	assign w49785 = w8993 ^ w8994;
	assign w46799 = w49785 ^ w995;
	assign w16064 = w46799 ^ w46797;
	assign w16139 = w16064 ^ w16154;
	assign w16130 = w16154 & w16139;
	assign w16039 = w16130 ^ w16131;
	assign w16026 = w16066 ^ w16064;
	assign w16142 = w16063 ^ w16026;
	assign w16138 = w46799 ^ w16065;
	assign w16134 = w16153 & w16138;
	assign w16068 = w16134 ^ w16064;
	assign w8969 = ~w9193;
	assign w8967 = w8969 ^ w49896;
	assign w8978 = w8969 ^ w9175;
	assign w49798 = w8967 ^ w8968;
	assign w46786 = w49798 ^ w1008;
	assign w16020 = w46786 ^ w46784;
	assign w49794 = w45352 ^ w8974;
	assign w46790 = w49794 ^ w1004;
	assign w8947 = w9171 ^ w9166;
	assign w8921 = w49892 ^ w8922;
	assign w9213 = w8920 ^ w8921;
	assign w49799 = w9213 ^ w9186;
	assign w46785 = w49799 ^ w1009;
	assign w49809 = w45359 ^ w8947;
	assign w15932 = w46784 ^ w46782;
	assign w15906 = w46785 ^ w46786;
	assign w9138 = w49884 ^ w49891;
	assign w8984 = w9197 ^ w9138;
	assign w49788 = w45346 ^ w8984;
	assign w46796 = w49788 ^ w998;
	assign w33088 = w46796 ^ w46790;
	assign w33165 = w33082 ^ w33088;
	assign w33168 = w46791 ^ w33088;
	assign w8946 = w9164 ^ w9160;
	assign w49810 = w45360 ^ w8946;
	assign w8945 = w9149 ^ w9138;
	assign w49811 = w49895 ^ w8945;
	assign w46773 = w49811 ^ w1021;
	assign w29953 = w46773 ^ w46778;
	assign w46775 = w49809 ^ w1019;
	assign w29866 = w46775 ^ w46773;
	assign w46774 = w49810 ^ w1020;
	assign w17091 = w46973 ^ w46979;
	assign w17072 = w17091 & w17076;
	assign w17006 = w17072 ^ w17002;
	assign w16980 = w17006 ^ w44081;
	assign w8966 = w49894 ^ w49888;
	assign w49801 = w8965 ^ w8966;
	assign w46783 = w49801 ^ w1011;
	assign w15891 = w15932 ^ w46783;
	assign w16040 = w46801 ^ w46802;
	assign w16086 = w16039 ^ w16040;
	assign w16085 = w16086 ^ w16068;
	assign w16129 = w16151 & w16142;
	assign w17005 = w17069 ^ w17003;
	assign w17064 = w16980 ^ w17005;
	assign w17011 = w17007 ^ w17005;
	assign w16979 = w17011 ^ w44084;
	assign w17016 = w46973 ^ w17011;
	assign w17066 = w17025 ^ w17016;
	assign w17022 = w46975 ^ w16979;
	assign w17024 = w16977 ^ w16978;
	assign w17023 = w17024 ^ w17006;
	assign w17065 = w17071 ^ w17023;
	assign w17062 = w17066 & w17065;
	assign w17057 = w17062 ^ w17022;
	assign w17056 = w17057 & w17058;
	assign w17054 = w17062 ^ w17056;
	assign w17053 = w17064 & w17054;
	assign w16975 = w17056 ^ w17020;
	assign w17055 = w17056 ^ w17064;
	assign w17041 = w17055 & w46980;
	assign w17032 = w17055 & w17087;
	assign w44083 = w17053 ^ w17071;
	assign w17045 = w44083 ^ w17023;
	assign w17034 = w17045 & w17086;
	assign w17043 = w17045 & w17082;
	assign w44086 = w17041 ^ w17043;
	assign w16974 = w17056 ^ w17073;
	assign w16025 = w16066 ^ w46799;
	assign w17012 = w46979 ^ w44083;
	assign w17052 = w17012 ^ w16975;
	assign w17042 = w17052 & w17081;
	assign w17033 = w17052 & w17083;
	assign w17061 = w17062 ^ w17064;
	assign w17060 = w17063 & w17061;
	assign w16968 = w17060 ^ w17016;
	assign w16971 = w17060 ^ w17072;
	assign w16967 = w16971 ^ w17007;
	assign w16966 = w46975 ^ w16967;
	assign w17059 = w17060 ^ w17022;
	assign w17038 = w17059 & w17078;
	assign w17029 = w17059 & w17085;
	assign w17051 = w17053 ^ w17061;
	assign w17050 = w17059 & w17051;
	assign w16973 = w17050 ^ w17074;
	assign w16965 = w17012 ^ w16973;
	assign w16972 = w17002 ^ w16965;
	assign w17044 = w16965 ^ w16966;
	assign w17027 = w17044 & w17092;
	assign w17036 = w17044 & w17077;
	assign w17015 = w17050 ^ w17025;
	assign w17046 = w17015 ^ w16968;
	assign w17031 = w17046 & w17091;
	assign w17040 = w17046 & w17076;
	assign w16998 = w17040 ^ w17031;
	assign w17049 = w17015 ^ w17017;
	assign w17039 = w17049 & w17088;
	assign w16997 = w17036 ^ w17039;
	assign w17030 = w17049 & w17084;
	assign w16982 = w17038 ^ w17039;
	assign w17000 = w17038 ^ w17030;
	assign w16994 = ~w16997;
	assign w16970 = w46973 ^ w16967;
	assign w44085 = w17039 ^ w17040;
	assign w17021 = w17036 ^ w44085;
	assign w16987 = w17032 ^ w17021;
	assign w16984 = ~w16987;
	assign w45777 = ~w33444;
	assign w9201 = w45346 ^ w45777;
	assign w8970 = w9201 ^ w9142;
	assign w49780 = w45777 ^ w8999;
	assign w8959 = w9201 ^ w9135;
	assign w49804 = w45354 ^ w8959;
	assign w46780 = w49804 ^ w1014;
	assign w29872 = w46780 ^ w46774;
	assign w29949 = w29866 ^ w29872;
	assign w29952 = w46775 ^ w29872;
	assign w8982 = w9201 ^ w9189;
	assign w8919 = w45354 ^ w45777;
	assign w9214 = w8918 ^ w8919;
	assign w49797 = w9214 ^ w9200;
	assign w46787 = w49797 ^ w1007;
	assign w15946 = w46787 ^ w46786;
	assign w15929 = w46787 ^ w46785;
	assign w15931 = w46786 ^ w15929;
	assign w16007 = w46782 ^ w15931;
	assign w46804 = w49780 ^ w990;
	assign w16070 = w46804 ^ w46798;
	assign w16140 = w16070 ^ w16065;
	assign w16150 = w46799 ^ w16070;
	assign w16146 = w46803 ^ w16150;
	assign w16133 = w16150 & w16146;
	assign w16127 = w16133 ^ w16085;
	assign w16147 = w16064 ^ w16070;
	assign w16145 = w16080 ^ w16147;
	assign w16132 = w16147 & w16140;
	assign w16143 = w46804 ^ w16144;
	assign w16136 = w16145 & w16143;
	assign w44042 = w16129 ^ w16132;
	assign w16082 = w16130 ^ w44042;
	assign w16038 = w16133 ^ w16082;
	assign w16120 = w46803 ^ w16038;
	assign w16042 = w16068 ^ w44042;
	assign w16004 = w46783 ^ w15931;
	assign w16149 = w46804 ^ w16025;
	assign w16135 = w46804 & w16149;
	assign w44041 = w16129 ^ w16135;
	assign w16079 = w44041 ^ w16064;
	assign w16126 = w16042 ^ w16067;
	assign w16041 = w16073 ^ w44041;
	assign w16084 = w46799 ^ w16041;
	assign w49796 = w45697 ^ w8970;
	assign w46788 = w49796 ^ w1006;
	assign w16015 = w46788 ^ w15891;
	assign w16001 = w46788 & w16015;
	assign w15936 = w46788 ^ w46782;
	assign w16016 = w46783 ^ w15936;
	assign w16012 = w46787 ^ w16016;
	assign w15999 = w16016 & w16012;
	assign w16006 = w15936 ^ w15931;
	assign w16087 = w16130 ^ w16136;
	assign w16125 = w16087 ^ w16079;
	assign w16128 = w16087 ^ w16078;
	assign w16124 = w16128 & w16127;
	assign w16123 = w16124 ^ w16126;
	assign w16119 = w16124 ^ w16084;
	assign w16118 = w16119 & w16120;
	assign w16036 = w16118 ^ w16135;
	assign w16037 = w16118 ^ w16082;
	assign w16117 = w16118 ^ w16126;
	assign w16103 = w16117 & w46804;
	assign w16094 = w16117 & w16149;
	assign w16031 = w16036 ^ w16132;
	assign w16122 = w16125 & w16123;
	assign w16030 = w16122 ^ w16078;
	assign w16121 = w16122 ^ w16084;
	assign w16100 = w16121 & w16140;
	assign w16091 = w16121 & w16147;
	assign w16033 = w16122 ^ w16134;
	assign w16029 = w16033 ^ w16069;
	assign w16028 = w46799 ^ w16029;
	assign w16032 = w46797 ^ w16029;
	assign w16109 = w16031 ^ w16032;
	assign w16099 = w16109 & w16141;
	assign w16090 = w16109 & w16152;
	assign w45897 = ~w9138;
	assign w8983 = w45897 ^ w45353;
	assign w8981 = w8982 ^ w8983;
	assign w49789 = ~w8981;
	assign w46795 = w49789 ^ w999;
	assign w33164 = w46795 ^ w33168;
	assign w33098 = w46795 ^ w46794;
	assign w33163 = w33098 ^ w33165;
	assign w33171 = w46789 ^ w46795;
	assign w33151 = w33168 & w33164;
	assign w8977 = w45897 ^ w49883;
	assign w49792 = w8976 ^ w8977;
	assign w46792 = w49792 ^ w1002;
	assign w33084 = w46792 ^ w46790;
	assign w33170 = w46792 ^ w46789;
	assign w33166 = w33170 ^ w33098;
	assign w33172 = w46794 ^ w46792;
	assign w33157 = w33082 ^ w33172;
	assign w33044 = w33084 ^ w33082;
	assign w33043 = w33084 ^ w46791;
	assign w33167 = w46796 ^ w33043;
	assign w33153 = w46796 & w33167;
	assign w33148 = w33172 & w33157;
	assign w8960 = w45897 ^ w49899;
	assign w49803 = w8960 ^ w8961;
	assign w46781 = w49803 ^ w1013;
	assign w15930 = w46783 ^ w46781;
	assign w16013 = w15930 ^ w15936;
	assign w16018 = w46784 ^ w46781;
	assign w16014 = w16018 ^ w15946;
	assign w16010 = w15929 ^ w16018;
	assign w16009 = w46788 ^ w16010;
	assign w15998 = w16013 & w16006;
	assign w16019 = w46781 ^ w46787;
	assign w16000 = w16019 & w16004;
	assign w15934 = w16000 ^ w15930;
	assign w15997 = w16018 & w16007;
	assign w15892 = w15932 ^ w15930;
	assign w16008 = w15929 ^ w15892;
	assign w16017 = w46781 ^ w46786;
	assign w15995 = w16017 & w16008;
	assign w16003 = w16010 & w16014;
	assign w8979 = w45897 ^ w49882;
	assign w49791 = w8978 ^ w8979;
	assign w44036 = w15995 ^ w16001;
	assign w44037 = w15995 ^ w15998;
	assign w15908 = w15934 ^ w44037;
	assign w15933 = w15997 ^ w15931;
	assign w15992 = w15908 ^ w15933;
	assign w16011 = w15946 ^ w16013;
	assign w16002 = w16011 & w16009;
	assign w46793 = w49791 ^ w1001;
	assign w33081 = w46795 ^ w46793;
	assign w33083 = w46794 ^ w33081;
	assign w33159 = w46790 ^ w33083;
	assign w33156 = w46791 ^ w33083;
	assign w33158 = w33088 ^ w33083;
	assign w33162 = w33081 ^ w33170;
	assign w33161 = w46796 ^ w33162;
	assign w33058 = w46793 ^ w46794;
	assign w33160 = w33081 ^ w33044;
	assign w33155 = w33162 & w33166;
	assign w33087 = w33155 ^ w33084;
	assign w33154 = w33163 & w33161;
	assign w33105 = w33148 ^ w33154;
	assign w33152 = w33171 & w33156;
	assign w33086 = w33152 ^ w33082;
	assign w33150 = w33165 & w33158;
	assign w33149 = w33170 & w33159;
	assign w33085 = w33149 ^ w33083;
	assign w33091 = w33087 ^ w33085;
	assign w33096 = w46789 ^ w33091;
	assign w33146 = w33105 ^ w33096;
	assign w33057 = w33148 ^ w33149;
	assign w33104 = w33057 ^ w33058;
	assign w33103 = w33104 ^ w33086;
	assign w33145 = w33151 ^ w33103;
	assign w33147 = w33169 & w33160;
	assign w33142 = w33146 & w33145;
	assign w44755 = w33147 ^ w33153;
	assign w33097 = w44755 ^ w33082;
	assign w33143 = w33105 ^ w33097;
	assign w33059 = w33091 ^ w44755;
	assign w33102 = w46791 ^ w33059;
	assign w33137 = w33142 ^ w33102;
	assign w44756 = w33147 ^ w33150;
	assign w33100 = w33148 ^ w44756;
	assign w33056 = w33151 ^ w33100;
	assign w33138 = w46795 ^ w33056;
	assign w33136 = w33137 & w33138;
	assign w33055 = w33136 ^ w33100;
	assign w33054 = w33136 ^ w33153;
	assign w33049 = w33054 ^ w33150;
	assign w33134 = w33142 ^ w33136;
	assign w33060 = w33086 ^ w44756;
	assign w33144 = w33060 ^ w33085;
	assign w33135 = w33136 ^ w33144;
	assign w33141 = w33142 ^ w33144;
	assign w33140 = w33143 & w33141;
	assign w33139 = w33140 ^ w33102;
	assign w33051 = w33140 ^ w33152;
	assign w33047 = w33051 ^ w33087;
	assign w33050 = w46789 ^ w33047;
	assign w33127 = w33049 ^ w33050;
	assign w33048 = w33140 ^ w33096;
	assign w33046 = w46791 ^ w33047;
	assign w33133 = w33144 & w33134;
	assign w33131 = w33133 ^ w33141;
	assign w33130 = w33139 & w33131;
	assign w33095 = w33130 ^ w33105;
	assign w33129 = w33095 ^ w33097;
	assign w33053 = w33130 ^ w33154;
	assign w33126 = w33095 ^ w33048;
	assign w33121 = w33135 & w46796;
	assign w33120 = w33126 & w33156;
	assign w33119 = w33129 & w33168;
	assign w33118 = w33139 & w33158;
	assign w33062 = w33118 ^ w33119;
	assign w33117 = w33127 & w33159;
	assign w33112 = w33135 & w33167;
	assign w33111 = w33126 & w33171;
	assign w33078 = w33120 ^ w33111;
	assign w33110 = w33129 & w33164;
	assign w33080 = w33118 ^ w33110;
	assign w33109 = w33139 & w33165;
	assign w33108 = w33127 & w33170;
	assign w44757 = w33119 ^ w33120;
	assign w44759 = w33133 ^ w33151;
	assign w33092 = w46795 ^ w44759;
	assign w33132 = w33092 ^ w33055;
	assign w33113 = w33132 & w33163;
	assign w33122 = w33132 & w33161;
	assign w33045 = w33092 ^ w33053;
	assign w33052 = w33082 ^ w33045;
	assign w33128 = w33049 ^ w33052;
	assign w33115 = w33128 & w33160;
	assign w33093 = w33111 ^ w33115;
	assign w33071 = ~w33093;
	assign w33070 = w33071 ^ w33109;
	assign w33124 = w33045 ^ w33046;
	assign w33107 = w33124 & w33172;
	assign w33106 = w33128 & w33169;
	assign w33072 = w33117 ^ w33106;
	assign w33068 = ~w33072;
	assign w43592 = w33107 ^ w33108;
	assign w33089 = w33113 ^ w43592;
	assign w33076 = w33080 ^ w43592;
	assign w33075 = w33071 ^ w33076;
	assign w33116 = w33124 & w33157;
	assign w33073 = w33116 ^ w33117;
	assign w33101 = w33116 ^ w44757;
	assign w33067 = w33112 ^ w33101;
	assign w33064 = ~w33067;
	assign w33061 = w33117 ^ w33101;
	assign w33077 = w33116 ^ w33119;
	assign w33074 = ~w33077;
	assign w33175 = w33074 ^ w33075;
	assign w33125 = w44759 ^ w33103;
	assign w33123 = w33125 & w33162;
	assign w33114 = w33125 & w33166;
	assign w33090 = w33114 ^ w33089;
	assign w33094 = w33122 ^ w33090;
	assign w33099 = w33123 ^ w33094;
	assign w50051 = w44757 ^ w33099;
	assign w33174 = w33099 ^ w33073;
	assign w33063 = w33121 ^ w33094;
	assign w50050 = w33062 ^ w33063;
	assign w50054 = w33090 ^ w33061;
	assign w50053 = ~w33174;
	assign w44758 = w33121 ^ w33123;
	assign w33079 = w44758 ^ w33076;
	assign w33176 = w33078 ^ w33079;
	assign w33066 = w33070 ^ w44758;
	assign w33069 = w33108 ^ w33066;
	assign w33173 = w33068 ^ w33069;
	assign w33065 = w33089 ^ w33066;
	assign w50049 = w33064 ^ w33065;
	assign w50052 = ~w33173;
	assign w15945 = w44036 ^ w15930;
	assign w16005 = w15930 ^ w16020;
	assign w15996 = w16020 & w16005;
	assign w15948 = w15996 ^ w44037;
	assign w15904 = w15999 ^ w15948;
	assign w15905 = w15996 ^ w15997;
	assign w15952 = w15905 ^ w15906;
	assign w15951 = w15952 ^ w15934;
	assign w15993 = w15999 ^ w15951;
	assign w15953 = w15996 ^ w16002;
	assign w15991 = w15953 ^ w15945;
	assign w15986 = w46787 ^ w15904;
	assign w45766 = ~w33176;
	assign w45773 = ~w33175;
	assign w16116 = w16124 ^ w16118;
	assign w16115 = w16126 & w16116;
	assign w16113 = w16115 ^ w16123;
	assign w16112 = w16121 & w16113;
	assign w16077 = w16112 ^ w16087;
	assign w16111 = w16077 ^ w16079;
	assign w16101 = w16111 & w16150;
	assign w16092 = w16111 & w16146;
	assign w16062 = w16100 ^ w16092;
	assign w16108 = w16077 ^ w16030;
	assign w16102 = w16108 & w16138;
	assign w16093 = w16108 & w16153;
	assign w16060 = w16102 ^ w16093;
	assign w16044 = w16100 ^ w16101;
	assign w16035 = w16112 ^ w16136;
	assign w44044 = w16101 ^ w16102;
	assign w44046 = w16115 ^ w16133;
	assign w16107 = w44046 ^ w16085;
	assign w16096 = w16107 & w16148;
	assign w16105 = w16107 & w16144;
	assign w44045 = w16103 ^ w16105;
	assign w16074 = w46803 ^ w44046;
	assign w16027 = w16074 ^ w16035;
	assign w16106 = w16027 ^ w16028;
	assign w16098 = w16106 & w16139;
	assign w16089 = w16106 & w16154;
	assign w16059 = w16098 ^ w16101;
	assign w16055 = w16098 ^ w16099;
	assign w16056 = ~w16059;
	assign w16034 = w16064 ^ w16027;
	assign w16110 = w16031 ^ w16034;
	assign w16088 = w16110 & w16151;
	assign w16054 = w16099 ^ w16088;
	assign w16050 = ~w16054;
	assign w16114 = w16074 ^ w16037;
	assign w16095 = w16114 & w16145;
	assign w16104 = w16114 & w16143;
	assign w16097 = w16110 & w16142;
	assign w16075 = w16093 ^ w16097;
	assign w16053 = ~w16075;
	assign w16052 = w16053 ^ w16091;
	assign w16048 = w16052 ^ w44045;
	assign w16051 = w16090 ^ w16048;
	assign w16155 = w16050 ^ w16051;
	assign w16083 = w16098 ^ w44044;
	assign w16049 = w16094 ^ w16083;
	assign w16046 = ~w16049;
	assign w16043 = w16099 ^ w16083;
	assign w44043 = w16089 ^ w16090;
	assign w16071 = w16095 ^ w44043;
	assign w16047 = w16071 ^ w16048;
	assign w16072 = w16096 ^ w16071;
	assign w16076 = w16104 ^ w16072;
	assign w16045 = w16103 ^ w16076;
	assign w50066 = w16044 ^ w16045;
	assign w50065 = w16046 ^ w16047;
	assign w16081 = w16105 ^ w16076;
	assign w50067 = w44044 ^ w16081;
	assign w16156 = w16081 ^ w16055;
	assign w16058 = w16062 ^ w44043;
	assign w16061 = w44045 ^ w16058;
	assign w16057 = w16053 ^ w16058;
	assign w16157 = w16056 ^ w16057;
	assign w16158 = w16060 ^ w16061;
	assign w50068 = w16072 ^ w16043;
	assign w45334 = ~w16155;
	assign w45335 = ~w16156;
	assign w9373 = w50068 ^ w45335;
	assign w45336 = ~w16157;
	assign w45337 = ~w16158;
	assign w15935 = w16003 ^ w15932;
	assign w15939 = w15935 ^ w15933;
	assign w15907 = w15939 ^ w44036;
	assign w15950 = w46783 ^ w15907;
	assign w15944 = w46781 ^ w15939;
	assign w15994 = w15953 ^ w15944;
	assign w15990 = w15994 & w15993;
	assign w15989 = w15990 ^ w15992;
	assign w15985 = w15990 ^ w15950;
	assign w15984 = w15985 & w15986;
	assign w15903 = w15984 ^ w15948;
	assign w15983 = w15984 ^ w15992;
	assign w15902 = w15984 ^ w16001;
	assign w15897 = w15902 ^ w15998;
	assign w15988 = w15991 & w15989;
	assign w15896 = w15988 ^ w15944;
	assign w15899 = w15988 ^ w16000;
	assign w15895 = w15899 ^ w15935;
	assign w15898 = w46781 ^ w15895;
	assign w15975 = w15897 ^ w15898;
	assign w15894 = w46783 ^ w15895;
	assign w15960 = w15983 & w16015;
	assign w15982 = w15990 ^ w15984;
	assign w15981 = w15992 & w15982;
	assign w15987 = w15988 ^ w15950;
	assign w15957 = w15987 & w16013;
	assign w15969 = w15983 & w46788;
	assign w15966 = w15987 & w16006;
	assign w44040 = w15981 ^ w15999;
	assign w15940 = w46787 ^ w44040;
	assign w15980 = w15940 ^ w15903;
	assign w15961 = w15980 & w16011;
	assign w15970 = w15980 & w16009;
	assign w15973 = w44040 ^ w15951;
	assign w15971 = w15973 & w16010;
	assign w44039 = w15969 ^ w15971;
	assign w15979 = w15981 ^ w15989;
	assign w15978 = w15987 & w15979;
	assign w15901 = w15978 ^ w16002;
	assign w15893 = w15940 ^ w15901;
	assign w15900 = w15930 ^ w15893;
	assign w15976 = w15897 ^ w15900;
	assign w15954 = w15976 & w16017;
	assign w15972 = w15893 ^ w15894;
	assign w15955 = w15972 & w16020;
	assign w15964 = w15972 & w16005;
	assign w15963 = w15976 & w16008;
	assign w15943 = w15978 ^ w15953;
	assign w15977 = w15943 ^ w15945;
	assign w15974 = w15943 ^ w15896;
	assign w15968 = w15974 & w16004;
	assign w15958 = w15977 & w16012;
	assign w15928 = w15966 ^ w15958;
	assign w15959 = w15974 & w16019;
	assign w15926 = w15968 ^ w15959;
	assign w15941 = w15959 ^ w15963;
	assign w15919 = ~w15941;
	assign w15918 = w15919 ^ w15957;
	assign w15914 = w15918 ^ w44039;
	assign w15967 = w15977 & w16016;
	assign w15910 = w15966 ^ w15967;
	assign w15925 = w15964 ^ w15967;
	assign w15922 = ~w15925;
	assign w44038 = w15967 ^ w15968;
	assign w15949 = w15964 ^ w44038;
	assign w15915 = w15960 ^ w15949;
	assign w15912 = ~w15915;
	assign w15956 = w15975 & w16018;
	assign w15917 = w15956 ^ w15914;
	assign w43543 = w15955 ^ w15956;
	assign w15937 = w15961 ^ w43543;
	assign w15913 = w15937 ^ w15914;
	assign w50110 = w15912 ^ w15913;
	assign w15924 = w15928 ^ w43543;
	assign w15927 = w44039 ^ w15924;
	assign w15923 = w15919 ^ w15924;
	assign w16023 = w15922 ^ w15923;
	assign w16024 = w15926 ^ w15927;
	assign w45332 = ~w16023;
	assign w45333 = ~w16024;
	assign w15965 = w15975 & w16007;
	assign w15920 = w15965 ^ w15954;
	assign w15916 = ~w15920;
	assign w15921 = w15964 ^ w15965;
	assign w15909 = w15965 ^ w15949;
	assign w16021 = w15916 ^ w15917;
	assign w45330 = ~w16021;
	assign w15962 = w15973 & w16014;
	assign w15938 = w15962 ^ w15937;
	assign w50113 = w15938 ^ w15909;
	assign w15942 = w15970 ^ w15938;
	assign w15947 = w15971 ^ w15942;
	assign w15911 = w15969 ^ w15942;
	assign w50111 = w15910 ^ w15911;
	assign w16022 = w15947 ^ w15921;
	assign w50112 = w44038 ^ w15947;
	assign w9286 = w50112 ^ w50111;
	assign w45331 = ~w16022;
	assign w9434 = w45331 ^ w45330;
	assign w16969 = w16974 ^ w17070;
	assign w17047 = w16969 ^ w16970;
	assign w17028 = w17047 & w17090;
	assign w17037 = w17047 & w17079;
	assign w16981 = w17037 ^ w17021;
	assign w17048 = w16969 ^ w16972;
	assign w17035 = w17048 & w17080;
	assign w17013 = w17031 ^ w17035;
	assign w17026 = w17048 & w17089;
	assign w16992 = w17037 ^ w17026;
	assign w16988 = ~w16992;
	assign w16991 = ~w17013;
	assign w16993 = w17036 ^ w17037;
	assign w16990 = w16991 ^ w17029;
	assign w16986 = w16990 ^ w44086;
	assign w16989 = w17028 ^ w16986;
	assign w17093 = w16988 ^ w16989;
	assign w44082 = w17027 ^ w17028;
	assign w16996 = w17000 ^ w44082;
	assign w16999 = w44086 ^ w16996;
	assign w17096 = w16998 ^ w16999;
	assign w16995 = w16991 ^ w16996;
	assign w17095 = w16994 ^ w16995;
	assign w17009 = w17033 ^ w44082;
	assign w16985 = w17009 ^ w16986;
	assign w17010 = w17034 ^ w17009;
	assign w49876 = w17010 ^ w16981;
	assign w17014 = w17042 ^ w17010;
	assign w16983 = w17041 ^ w17014;
	assign w17019 = w17043 ^ w17014;
	assign w9144 = w49872 ^ w49876;
	assign w9136 = w49876 ^ w49880;
	assign w49873 = w16984 ^ w16985;
	assign w17094 = w17019 ^ w16993;
	assign w49874 = w16982 ^ w16983;
	assign w49875 = w44085 ^ w17019;
	assign w9157 = w49875 ^ w49879;
	assign w49752 = w9223 ^ w9157;
	assign w9162 = w49874 ^ w49878;
	assign w49751 = w9224 ^ w9162;
	assign w46832 = w49752 ^ w1026;
	assign w46833 = w49751 ^ w1025;
	assign w9167 = w49873 ^ w49877;
	assign w9050 = w9167 ^ w45524;
	assign w49750 = w9050 ^ w9051;
	assign w46834 = w49750 ^ w1024;
	assign w16288 = w46834 ^ w46832;
	assign w16174 = w46833 ^ w46834;
	assign w9034 = w9025 ^ w9162;
	assign w9045 = w9155 ^ w9136;
	assign w49755 = w49872 ^ w9045;
	assign w46829 = w49755 ^ w1029;
	assign w16285 = w46829 ^ w46834;
	assign w16286 = w46832 ^ w46829;
	assign w9027 = w9136 ^ w45771;
	assign w9031 = w9033 ^ w9157;
	assign w9006 = ~w49875;
	assign w9026 = w9177 ^ w9144;
	assign w49764 = w45525 ^ w9026;
	assign w9012 = w9136 ^ w49874;
	assign w9016 = w9177 ^ w9136;
	assign w49763 = w9027 ^ w9028;
	assign w9021 = w9006 ^ w49871;
	assign w49769 = w9020 ^ w9021;
	assign w46815 = w49769 ^ w1043;
	assign w9004 = w9007 ^ w9162;
	assign w9005 = w9136 ^ w9006;
	assign w49776 = w9004 ^ w9005;
	assign w46808 = w49776 ^ w1050;
	assign w9003 = w9161 ^ w9157;
	assign w9036 = w9176 ^ w9167;
	assign w49758 = w49864 ^ w9036;
	assign w8906 = w49873 ^ w49869;
	assign w8909 = ~w9144;
	assign w8907 = w8909 ^ w49879;
	assign w8908 = w49874 ^ w8896;
	assign w9218 = w8907 ^ w8908;
	assign w49768 = w9218 ^ w9165;
	assign w8905 = w9144 ^ w49878;
	assign w9219 = w8905 ^ w8906;
	assign w49767 = w9219 ^ w9169;
	assign w46817 = w49767 ^ w1041;
	assign w8903 = w9144 ^ w45524;
	assign w46816 = w49768 ^ w1042;
	assign w46826 = w49758 ^ w1032;
	assign w46820 = w49764 ^ w1038;
	assign w46821 = w49763 ^ w1037;
	assign w9011 = w9169 ^ w9167;
	assign w49775 = w9011 ^ w9012;
	assign w46809 = w49775 ^ w1049;
	assign w45358 = ~w17096;
	assign w9174 = w45358 ^ w45525;
	assign w9052 = w9174 ^ w9146;
	assign w49748 = w45772 ^ w9052;
	assign w46836 = w49748 ^ w1022;
	assign w49772 = w45358 ^ w9016;
	assign w46812 = w49772 ^ w1046;
	assign w9040 = w9174 ^ w9137;
	assign w49756 = w45350 ^ w9040;
	assign w46828 = w49756 ^ w1030;
	assign w9014 = w9176 ^ w9174;
	assign w8904 = w45358 ^ w45772;
	assign w9220 = w8903 ^ w8904;
	assign w49765 = w9220 ^ w9176;
	assign w46819 = w49765 ^ w1039;
	assign w45363 = ~w17093;
	assign w9152 = w45363 ^ w45522;
	assign w49777 = w45363 ^ w9003;
	assign w46807 = w49777 ^ w1051;
	assign w9030 = w9165 ^ w9152;
	assign w49761 = w45355 ^ w9030;
	assign w46823 = w49761 ^ w1035;
	assign w11642 = w46823 ^ w46821;
	assign w9018 = w9155 ^ w45363;
	assign w49770 = w9018 ^ w9019;
	assign w46814 = w49770 ^ w1044;
	assign w26920 = w46816 ^ w46814;
	assign w26924 = w46820 ^ w46814;
	assign w27004 = w46815 ^ w26924;
	assign w27000 = w46819 ^ w27004;
	assign w26987 = w27004 & w27000;
	assign w26879 = w26920 ^ w46815;
	assign w27003 = w46820 ^ w26879;
	assign w9048 = w9152 ^ w49879;
	assign w49753 = w9048 ^ w9049;
	assign w46831 = w49753 ^ w1027;
	assign w16198 = w46831 ^ w46829;
	assign w16273 = w16198 ^ w16288;
	assign w16264 = w16288 & w16273;
	assign w26989 = w46820 & w27003;
	assign w45364 = ~w17094;
	assign w9001 = w49876 ^ w45364;
	assign w49762 = w45364 ^ w9029;
	assign w49779 = w9000 ^ w9001;
	assign w46805 = w49779 ^ w1053;
	assign w30000 = w46807 ^ w46805;
	assign w30088 = w46808 ^ w46805;
	assign w46822 = w49762 ^ w1036;
	assign w11648 = w46828 ^ w46822;
	assign w11725 = w11642 ^ w11648;
	assign w11728 = w46823 ^ w11648;
	assign w9154 = w45771 ^ w45364;
	assign w9046 = w9154 ^ w45523;
	assign w49754 = w9046 ^ w9047;
	assign w46830 = w49754 ^ w1028;
	assign w16204 = w46836 ^ w46830;
	assign w16284 = w46831 ^ w16204;
	assign w16200 = w46832 ^ w46830;
	assign w16160 = w16200 ^ w16198;
	assign w16159 = w16200 ^ w46831;
	assign w9002 = w9154 ^ w9152;
	assign w49778 = w45356 ^ w9002;
	assign w46806 = w49778 ^ w1052;
	assign w30002 = w46808 ^ w46806;
	assign w30006 = w46812 ^ w46806;
	assign w30083 = w30000 ^ w30006;
	assign w30086 = w46807 ^ w30006;
	assign w29962 = w30002 ^ w30000;
	assign w29961 = w30002 ^ w46807;
	assign w30085 = w46812 ^ w29961;
	assign w30071 = w46812 & w30085;
	assign w16281 = w16198 ^ w16204;
	assign w9017 = w9154 ^ w9137;
	assign w49771 = w49880 ^ w9017;
	assign w46813 = w49771 ^ w1045;
	assign w27006 = w46816 ^ w46813;
	assign w27007 = w46813 ^ w46819;
	assign w26918 = w46815 ^ w46813;
	assign w27001 = w26918 ^ w26924;
	assign w26880 = w26920 ^ w26918;
	assign w16283 = w46836 ^ w16159;
	assign w16269 = w46836 & w16283;
	assign w45365 = ~w17095;
	assign w9170 = w45365 ^ w45524;
	assign w49749 = w9225 ^ w9170;
	assign w46835 = w49749 ^ w1023;
	assign w16197 = w46835 ^ w46833;
	assign w16280 = w46835 ^ w16284;
	assign w16278 = w16197 ^ w16286;
	assign w16214 = w46835 ^ w46834;
	assign w16279 = w16214 ^ w16281;
	assign w16199 = w46834 ^ w16197;
	assign w16274 = w16204 ^ w16199;
	assign w16266 = w16281 & w16274;
	assign w16275 = w46830 ^ w16199;
	assign w16265 = w16286 & w16275;
	assign w16272 = w46831 ^ w16199;
	assign w16287 = w46829 ^ w46835;
	assign w16201 = w16265 ^ w16199;
	assign w16268 = w16287 & w16272;
	assign w16202 = w16268 ^ w16198;
	assign w16173 = w16264 ^ w16265;
	assign w16220 = w16173 ^ w16174;
	assign w16219 = w16220 ^ w16202;
	assign w16267 = w16284 & w16280;
	assign w16261 = w16267 ^ w16219;
	assign w9015 = w9136 ^ w45365;
	assign w9038 = w9177 ^ w9170;
	assign w9024 = w45365 ^ w33309;
	assign w49766 = w9023 ^ w9024;
	assign w46818 = w49766 ^ w1040;
	assign w26894 = w46817 ^ w46818;
	assign w26934 = w46819 ^ w46818;
	assign w27008 = w46818 ^ w46816;
	assign w27002 = w27006 ^ w26934;
	assign w49773 = w9014 ^ w9015;
	assign w46811 = w49773 ^ w1047;
	assign w29999 = w46811 ^ w46809;
	assign w30082 = w46811 ^ w30086;
	assign w30080 = w29999 ^ w30088;
	assign w30079 = w46812 ^ w30080;
	assign w30078 = w29999 ^ w29962;
	assign w30089 = w46805 ^ w46811;
	assign w30069 = w30086 & w30082;
	assign w9013 = w9172 ^ w9170;
	assign w49774 = w49873 ^ w9013;
	assign w46810 = w49774 ^ w1048;
	assign w30001 = w46810 ^ w29999;
	assign w30077 = w46806 ^ w30001;
	assign w30074 = w46807 ^ w30001;
	assign w30076 = w30006 ^ w30001;
	assign w30016 = w46811 ^ w46810;
	assign w30081 = w30016 ^ w30083;
	assign w30084 = w30088 ^ w30016;
	assign w30090 = w46810 ^ w46808;
	assign w30075 = w30000 ^ w30090;
	assign w29976 = w46809 ^ w46810;
	assign w30087 = w46805 ^ w46810;
	assign w30073 = w30080 & w30084;
	assign w30005 = w30073 ^ w30002;
	assign w30072 = w30081 & w30079;
	assign w30070 = w30089 & w30074;
	assign w30004 = w30070 ^ w30000;
	assign w30068 = w30083 & w30076;
	assign w30067 = w30088 & w30077;
	assign w30003 = w30067 ^ w30001;
	assign w30009 = w30005 ^ w30003;
	assign w30014 = w46805 ^ w30009;
	assign w30066 = w30090 & w30075;
	assign w30023 = w30066 ^ w30072;
	assign w30064 = w30023 ^ w30014;
	assign w29975 = w30066 ^ w30067;
	assign w30022 = w29975 ^ w29976;
	assign w30021 = w30022 ^ w30004;
	assign w30063 = w30069 ^ w30021;
	assign w30065 = w30087 & w30078;
	assign w30060 = w30064 & w30063;
	assign w26999 = w26934 ^ w27001;
	assign w27005 = w46813 ^ w46818;
	assign w16282 = w16286 ^ w16214;
	assign w16276 = w16197 ^ w16160;
	assign w16263 = w16285 & w16276;
	assign w44047 = w16263 ^ w16266;
	assign w16176 = w16202 ^ w44047;
	assign w16260 = w16176 ^ w16201;
	assign w44050 = w16263 ^ w16269;
	assign w16213 = w44050 ^ w16198;
	assign w16216 = w16264 ^ w44047;
	assign w16172 = w16267 ^ w16216;
	assign w16254 = w46835 ^ w16172;
	assign w16271 = w16278 & w16282;
	assign w16203 = w16271 ^ w16200;
	assign w16207 = w16203 ^ w16201;
	assign w16212 = w46829 ^ w16207;
	assign w16175 = w16207 ^ w44050;
	assign w16218 = w46831 ^ w16175;
	assign w44626 = w30065 ^ w30068;
	assign w29978 = w30004 ^ w44626;
	assign w30062 = w29978 ^ w30003;
	assign w30059 = w30060 ^ w30062;
	assign w30018 = w30066 ^ w44626;
	assign w29974 = w30069 ^ w30018;
	assign w30056 = w46811 ^ w29974;
	assign w44629 = w30065 ^ w30071;
	assign w29977 = w30009 ^ w44629;
	assign w30020 = w46807 ^ w29977;
	assign w30055 = w30060 ^ w30020;
	assign w30054 = w30055 & w30056;
	assign w30052 = w30060 ^ w30054;
	assign w29973 = w30054 ^ w30018;
	assign w29972 = w30054 ^ w30071;
	assign w29967 = w29972 ^ w30068;
	assign w30051 = w30062 & w30052;
	assign w30049 = w30051 ^ w30059;
	assign w44628 = w30051 ^ w30069;
	assign w30043 = w44628 ^ w30021;
	assign w30032 = w30043 & w30084;
	assign w30041 = w30043 & w30080;
	assign w30010 = w46811 ^ w44628;
	assign w30050 = w30010 ^ w29973;
	assign w30040 = w30050 & w30079;
	assign w30031 = w30050 & w30081;
	assign w30053 = w30054 ^ w30062;
	assign w30039 = w30053 & w46812;
	assign w30030 = w30053 & w30085;
	assign w30015 = w44629 ^ w30000;
	assign w30061 = w30023 ^ w30015;
	assign w30058 = w30061 & w30059;
	assign w30057 = w30058 ^ w30020;
	assign w29969 = w30058 ^ w30070;
	assign w29965 = w29969 ^ w30005;
	assign w29968 = w46805 ^ w29965;
	assign w30045 = w29967 ^ w29968;
	assign w29966 = w30058 ^ w30014;
	assign w29964 = w46807 ^ w29965;
	assign w30048 = w30057 & w30049;
	assign w30013 = w30048 ^ w30023;
	assign w30047 = w30013 ^ w30015;
	assign w29971 = w30048 ^ w30072;
	assign w29963 = w30010 ^ w29971;
	assign w29970 = w30000 ^ w29963;
	assign w30046 = w29967 ^ w29970;
	assign w30044 = w30013 ^ w29966;
	assign w30042 = w29963 ^ w29964;
	assign w30038 = w30044 & w30074;
	assign w30037 = w30047 & w30086;
	assign w30036 = w30057 & w30076;
	assign w29980 = w30036 ^ w30037;
	assign w30035 = w30045 & w30077;
	assign w30034 = w30042 & w30075;
	assign w29995 = w30034 ^ w30037;
	assign w29992 = ~w29995;
	assign w29991 = w30034 ^ w30035;
	assign w30033 = w30046 & w30078;
	assign w30029 = w30044 & w30089;
	assign w30011 = w30029 ^ w30033;
	assign w29996 = w30038 ^ w30029;
	assign w29989 = ~w30011;
	assign w30028 = w30047 & w30082;
	assign w29998 = w30036 ^ w30028;
	assign w30027 = w30057 & w30083;
	assign w29988 = w29989 ^ w30027;
	assign w30026 = w30045 & w30088;
	assign w30025 = w30042 & w30090;
	assign w30024 = w30046 & w30087;
	assign w29990 = w30035 ^ w30024;
	assign w29986 = ~w29990;
	assign w44627 = w30025 ^ w30026;
	assign w30007 = w30031 ^ w44627;
	assign w30008 = w30032 ^ w30007;
	assign w30012 = w30040 ^ w30008;
	assign w29981 = w30039 ^ w30012;
	assign w50079 = w29980 ^ w29981;
	assign w30017 = w30041 ^ w30012;
	assign w30092 = w30017 ^ w29991;
	assign w29994 = w29998 ^ w44627;
	assign w29993 = w29989 ^ w29994;
	assign w30093 = w29992 ^ w29993;
	assign w44630 = w30037 ^ w30038;
	assign w50080 = w44630 ^ w30017;
	assign w30019 = w30034 ^ w44630;
	assign w29985 = w30030 ^ w30019;
	assign w29982 = ~w29985;
	assign w29979 = w30035 ^ w30019;
	assign w50081 = w30008 ^ w29979;
	assign w9491 = w50068 ^ w50081;
	assign w9238 = ~w9491;
	assign w44631 = w30039 ^ w30041;
	assign w29997 = w44631 ^ w29994;
	assign w30094 = w29996 ^ w29997;
	assign w29984 = w29988 ^ w44631;
	assign w29987 = w30026 ^ w29984;
	assign w30091 = w29986 ^ w29987;
	assign w29983 = w30007 ^ w29984;
	assign w50078 = w29982 ^ w29983;
	assign w9239 = w9238 ^ w50078;
	assign w26993 = w26918 ^ w27008;
	assign w26984 = w27008 & w26993;
	assign w16277 = w46836 ^ w16278;
	assign w16270 = w16279 & w16277;
	assign w16221 = w16264 ^ w16270;
	assign w16259 = w16221 ^ w16213;
	assign w16262 = w16221 ^ w16212;
	assign w16258 = w16262 & w16261;
	assign w16253 = w16258 ^ w16218;
	assign w16257 = w16258 ^ w16260;
	assign w16256 = w16259 & w16257;
	assign w16167 = w16256 ^ w16268;
	assign w16163 = w16167 ^ w16203;
	assign w16252 = w16253 & w16254;
	assign w16170 = w16252 ^ w16269;
	assign w16165 = w16170 ^ w16266;
	assign w16250 = w16258 ^ w16252;
	assign w16249 = w16260 & w16250;
	assign w16255 = w16256 ^ w16218;
	assign w16234 = w16255 & w16274;
	assign w16251 = w16252 ^ w16260;
	assign w16237 = w16251 & w46836;
	assign w16171 = w16252 ^ w16216;
	assign w16247 = w16249 ^ w16257;
	assign w16246 = w16255 & w16247;
	assign w16211 = w16246 ^ w16221;
	assign w16245 = w16211 ^ w16213;
	assign w16169 = w16246 ^ w16270;
	assign w16235 = w16245 & w16284;
	assign w16228 = w16251 & w16283;
	assign w16164 = w16256 ^ w16212;
	assign w16242 = w16211 ^ w16164;
	assign w16227 = w16242 & w16287;
	assign w16236 = w16242 & w16272;
	assign w16194 = w16236 ^ w16227;
	assign w44049 = w16249 ^ w16267;
	assign w16241 = w44049 ^ w16219;
	assign w16230 = w16241 & w16282;
	assign w16239 = w16241 & w16278;
	assign w16208 = w46835 ^ w44049;
	assign w16161 = w16208 ^ w16169;
	assign w16248 = w16208 ^ w16171;
	assign w16238 = w16248 & w16277;
	assign w44051 = w16235 ^ w16236;
	assign w44052 = w16237 ^ w16239;
	assign w16225 = w16255 & w16281;
	assign w16226 = w16245 & w16280;
	assign w16196 = w16234 ^ w16226;
	assign w16229 = w16248 & w16279;
	assign w9242 = w9491 ^ w50079;
	assign w45686 = ~w30091;
	assign w9392 = w45686 ^ w45334;
	assign w45687 = ~w30092;
	assign w9500 = w45335 ^ w45687;
	assign w45688 = ~w30093;
	assign w45689 = ~w30094;
	assign w9236 = w9238 ^ w45689;
	assign w16178 = w16234 ^ w16235;
	assign w16166 = w46829 ^ w16163;
	assign w16243 = w16165 ^ w16166;
	assign w16233 = w16243 & w16275;
	assign w16224 = w16243 & w16286;
	assign w16162 = w46831 ^ w16163;
	assign w16240 = w16161 ^ w16162;
	assign w16232 = w16240 & w16273;
	assign w16189 = w16232 ^ w16233;
	assign w16217 = w16232 ^ w44051;
	assign w16183 = w16228 ^ w16217;
	assign w16180 = ~w16183;
	assign w16193 = w16232 ^ w16235;
	assign w16190 = ~w16193;
	assign w16223 = w16240 & w16288;
	assign w44048 = w16223 ^ w16224;
	assign w16205 = w16229 ^ w44048;
	assign w16206 = w16230 ^ w16205;
	assign w16210 = w16238 ^ w16206;
	assign w16215 = w16239 ^ w16210;
	assign w16290 = w16215 ^ w16189;
	assign w50047 = w44051 ^ w16215;
	assign w9540 = w50047 ^ w50051;
	assign w16192 = w16196 ^ w44048;
	assign w16195 = w44052 ^ w16192;
	assign w16292 = w16194 ^ w16195;
	assign w45339 = ~w16290;
	assign w9535 = w45339 ^ w50053;
	assign w45341 = ~w16292;
	assign w16177 = w16233 ^ w16217;
	assign w16179 = w16237 ^ w16210;
	assign w50046 = w16178 ^ w16179;
	assign w9549 = w50046 ^ w50050;
	assign w9431 = ~w9549;
	assign w50048 = w16206 ^ w16177;
	assign w9485 = w50048 ^ w50054;
	assign w9275 = w9485 ^ w50046;
	assign w11729 = w46821 ^ w46826;
	assign w26917 = w46819 ^ w46817;
	assign w26998 = w26917 ^ w27006;
	assign w26919 = w46818 ^ w26917;
	assign w26994 = w26924 ^ w26919;
	assign w26992 = w46815 ^ w26919;
	assign w26986 = w27001 & w26994;
	assign w26991 = w26998 & w27002;
	assign w26995 = w46814 ^ w26919;
	assign w26985 = w27006 & w26995;
	assign w26893 = w26984 ^ w26985;
	assign w26921 = w26985 ^ w26919;
	assign w26997 = w46820 ^ w26998;
	assign w26923 = w26991 ^ w26920;
	assign w26996 = w26917 ^ w26880;
	assign w26983 = w27005 & w26996;
	assign w44496 = w26983 ^ w26989;
	assign w26933 = w44496 ^ w26918;
	assign w44497 = w26983 ^ w26986;
	assign w26936 = w26984 ^ w44497;
	assign w26927 = w26923 ^ w26921;
	assign w26932 = w46813 ^ w26927;
	assign w26895 = w26927 ^ w44496;
	assign w26940 = w26893 ^ w26894;
	assign w26990 = w26999 & w26997;
	assign w26941 = w26984 ^ w26990;
	assign w26982 = w26941 ^ w26932;
	assign w26979 = w26941 ^ w26933;
	assign w26938 = w46815 ^ w26895;
	assign w26892 = w26987 ^ w26936;
	assign w26974 = w46819 ^ w26892;
	assign w26988 = w27007 & w26992;
	assign w26922 = w26988 ^ w26918;
	assign w26939 = w26940 ^ w26922;
	assign w26981 = w26987 ^ w26939;
	assign w26978 = w26982 & w26981;
	assign w26973 = w26978 ^ w26938;
	assign w26896 = w26922 ^ w44497;
	assign w26980 = w26896 ^ w26921;
	assign w26977 = w26978 ^ w26980;
	assign w26976 = w26979 & w26977;
	assign w26884 = w26976 ^ w26932;
	assign w26887 = w26976 ^ w26988;
	assign w26883 = w26887 ^ w26923;
	assign w26882 = w46815 ^ w26883;
	assign w26886 = w46813 ^ w26883;
	assign w26975 = w26976 ^ w26938;
	assign w26945 = w26975 & w27001;
	assign w26954 = w26975 & w26994;
	assign w26972 = w26973 & w26974;
	assign w26890 = w26972 ^ w26989;
	assign w26885 = w26890 ^ w26986;
	assign w26963 = w26885 ^ w26886;
	assign w26953 = w26963 & w26995;
	assign w26944 = w26963 & w27006;
	assign w26891 = w26972 ^ w26936;
	assign w26971 = w26972 ^ w26980;
	assign w26957 = w26971 & w46820;
	assign w26948 = w26971 & w27003;
	assign w26970 = w26978 ^ w26972;
	assign w26969 = w26980 & w26970;
	assign w26967 = w26969 ^ w26977;
	assign w26966 = w26975 & w26967;
	assign w26889 = w26966 ^ w26990;
	assign w26931 = w26966 ^ w26941;
	assign w26962 = w26931 ^ w26884;
	assign w26947 = w26962 & w27007;
	assign w26965 = w26931 ^ w26933;
	assign w26946 = w26965 & w27000;
	assign w26916 = w26954 ^ w26946;
	assign w26955 = w26965 & w27004;
	assign w26898 = w26954 ^ w26955;
	assign w26956 = w26962 & w26992;
	assign w26914 = w26956 ^ w26947;
	assign w44498 = w26955 ^ w26956;
	assign w44500 = w26969 ^ w26987;
	assign w26928 = w46819 ^ w44500;
	assign w26968 = w26928 ^ w26891;
	assign w26958 = w26968 & w26997;
	assign w26881 = w26928 ^ w26889;
	assign w26960 = w26881 ^ w26882;
	assign w26943 = w26960 & w27008;
	assign w43575 = w26943 ^ w26944;
	assign w26912 = w26916 ^ w43575;
	assign w26952 = w26960 & w26993;
	assign w26937 = w26952 ^ w44498;
	assign w26903 = w26948 ^ w26937;
	assign w26900 = ~w26903;
	assign w26913 = w26952 ^ w26955;
	assign w26909 = w26952 ^ w26953;
	assign w26897 = w26953 ^ w26937;
	assign w26910 = ~w26913;
	assign w26949 = w26968 & w26999;
	assign w26925 = w26949 ^ w43575;
	assign w26961 = w44500 ^ w26939;
	assign w26950 = w26961 & w27002;
	assign w26926 = w26950 ^ w26925;
	assign w26930 = w26958 ^ w26926;
	assign w26899 = w26957 ^ w26930;
	assign w50094 = w26898 ^ w26899;
	assign w50096 = w26926 ^ w26897;
	assign w26888 = w26918 ^ w26881;
	assign w26964 = w26885 ^ w26888;
	assign w26942 = w26964 & w27005;
	assign w26908 = w26953 ^ w26942;
	assign w26951 = w26964 & w26996;
	assign w26929 = w26947 ^ w26951;
	assign w26907 = ~w26929;
	assign w26906 = w26907 ^ w26945;
	assign w26911 = w26907 ^ w26912;
	assign w27011 = w26910 ^ w26911;
	assign w26904 = ~w26908;
	assign w45598 = ~w27011;
	assign w26959 = w26961 & w26998;
	assign w26935 = w26959 ^ w26930;
	assign w50095 = w44498 ^ w26935;
	assign w27010 = w26935 ^ w26909;
	assign w44499 = w26957 ^ w26959;
	assign w26915 = w44499 ^ w26912;
	assign w27012 = w26914 ^ w26915;
	assign w26902 = w26906 ^ w44499;
	assign w26901 = w26925 ^ w26902;
	assign w26905 = w26944 ^ w26902;
	assign w27009 = w26904 ^ w26905;
	assign w50093 = w26900 ^ w26901;
	assign w45599 = ~w27012;
	assign w45604 = ~w27009;
	assign w45605 = ~w27010;
	assign w16168 = w16198 ^ w16161;
	assign w16244 = w16165 ^ w16168;
	assign w16231 = w16244 & w16276;
	assign w16209 = w16227 ^ w16231;
	assign w16187 = ~w16209;
	assign w16186 = w16187 ^ w16225;
	assign w16182 = w16186 ^ w44052;
	assign w16181 = w16205 ^ w16182;
	assign w16222 = w16244 & w16285;
	assign w16188 = w16233 ^ w16222;
	assign w16184 = ~w16188;
	assign w16191 = w16187 ^ w16192;
	assign w16291 = w16190 ^ w16191;
	assign w50045 = w16180 ^ w16181;
	assign w9276 = w50045 ^ w50049;
	assign w9554 = w9275 ^ w9276;
	assign w45340 = ~w16291;
	assign w16185 = w16224 ^ w16182;
	assign w16289 = w16184 ^ w16185;
	assign w45338 = ~w16289;
	assign w9537 = w45338 ^ w50052;
	assign w45937 = ~w8795;
	assign w8590 = w45937 ^ w49658;
	assign w8863 = w8590 ^ w8591;
	assign w8714 = w45937 ^ w49656;
	assign w49543 = w8713 ^ w8714;
	assign w8627 = w45937 ^ w45389;
	assign w49522 = w8627 ^ w8628;
	assign w46989 = w49522 ^ w934;
	assign w17136 = w46991 ^ w46989;
	assign w17211 = w17136 ^ w17226;
	assign w17219 = w17136 ^ w17142;
	assign w17217 = w17152 ^ w17219;
	assign w17224 = w46992 ^ w46989;
	assign w17220 = w17224 ^ w17152;
	assign w17216 = w17135 ^ w17224;
	assign w17215 = w46996 ^ w17216;
	assign w17223 = w46989 ^ w46994;
	assign w17225 = w46989 ^ w46995;
	assign w17098 = w17138 ^ w17136;
	assign w17214 = w17135 ^ w17098;
	assign w17208 = w17217 & w17215;
	assign w17209 = w17216 & w17220;
	assign w17141 = w17209 ^ w17138;
	assign w17206 = w17225 & w17210;
	assign w17140 = w17206 ^ w17136;
	assign w17204 = w17219 & w17212;
	assign w17203 = w17224 & w17213;
	assign w17139 = w17203 ^ w17137;
	assign w17145 = w17141 ^ w17139;
	assign w17150 = w46989 ^ w17145;
	assign w17202 = w17226 & w17211;
	assign w17111 = w17202 ^ w17203;
	assign w17158 = w17111 ^ w17112;
	assign w17159 = w17202 ^ w17208;
	assign w17200 = w17159 ^ w17150;
	assign w17157 = w17158 ^ w17140;
	assign w17199 = w17205 ^ w17157;
	assign w17196 = w17200 & w17199;
	assign w46968 = w49543 ^ w955;
	assign w30404 = w46968 ^ w46966;
	assign w30490 = w46968 ^ w46965;
	assign w30486 = w30490 ^ w30418;
	assign w30492 = w46970 ^ w46968;
	assign w30477 = w30402 ^ w30492;
	assign w30364 = w30404 ^ w30402;
	assign w30363 = w30404 ^ w46967;
	assign w30487 = w46972 ^ w30363;
	assign w30473 = w46972 & w30487;
	assign w30468 = w30492 & w30477;
	assign w49542 = w8863 ^ w8860;
	assign w46969 = w49542 ^ w954;
	assign w30401 = w46971 ^ w46969;
	assign w30403 = w46970 ^ w30401;
	assign w30479 = w46966 ^ w30403;
	assign w30476 = w46967 ^ w30403;
	assign w30478 = w30408 ^ w30403;
	assign w30482 = w30401 ^ w30490;
	assign w30481 = w46972 ^ w30482;
	assign w30378 = w46969 ^ w46970;
	assign w30480 = w30401 ^ w30364;
	assign w30475 = w30482 & w30486;
	assign w30407 = w30475 ^ w30404;
	assign w30474 = w30483 & w30481;
	assign w30425 = w30468 ^ w30474;
	assign w30472 = w30491 & w30476;
	assign w30406 = w30472 ^ w30402;
	assign w30470 = w30485 & w30478;
	assign w30469 = w30490 & w30479;
	assign w30405 = w30469 ^ w30403;
	assign w30411 = w30407 ^ w30405;
	assign w30416 = w46965 ^ w30411;
	assign w30466 = w30425 ^ w30416;
	assign w30377 = w30468 ^ w30469;
	assign w30424 = w30377 ^ w30378;
	assign w30423 = w30424 ^ w30406;
	assign w30465 = w30471 ^ w30423;
	assign w30467 = w30489 & w30480;
	assign w30462 = w30466 & w30465;
	assign w44643 = w30467 ^ w30470;
	assign w30380 = w30406 ^ w44643;
	assign w30464 = w30380 ^ w30405;
	assign w30461 = w30462 ^ w30464;
	assign w30420 = w30468 ^ w44643;
	assign w30376 = w30471 ^ w30420;
	assign w30458 = w46971 ^ w30376;
	assign w44646 = w30467 ^ w30473;
	assign w30379 = w30411 ^ w44646;
	assign w30422 = w46967 ^ w30379;
	assign w30457 = w30462 ^ w30422;
	assign w30456 = w30457 & w30458;
	assign w30454 = w30462 ^ w30456;
	assign w30375 = w30456 ^ w30420;
	assign w30374 = w30456 ^ w30473;
	assign w30369 = w30374 ^ w30470;
	assign w30453 = w30464 & w30454;
	assign w30451 = w30453 ^ w30461;
	assign w44645 = w30453 ^ w30471;
	assign w30445 = w44645 ^ w30423;
	assign w30434 = w30445 & w30486;
	assign w30443 = w30445 & w30482;
	assign w30412 = w46971 ^ w44645;
	assign w30452 = w30412 ^ w30375;
	assign w30442 = w30452 & w30481;
	assign w30433 = w30452 & w30483;
	assign w30455 = w30456 ^ w30464;
	assign w30441 = w30455 & w46972;
	assign w30432 = w30455 & w30487;
	assign w30417 = w44646 ^ w30402;
	assign w30463 = w30425 ^ w30417;
	assign w30460 = w30463 & w30461;
	assign w30459 = w30460 ^ w30422;
	assign w30371 = w30460 ^ w30472;
	assign w30367 = w30371 ^ w30407;
	assign w30370 = w46965 ^ w30367;
	assign w30447 = w30369 ^ w30370;
	assign w30368 = w30460 ^ w30416;
	assign w30366 = w46967 ^ w30367;
	assign w30450 = w30459 & w30451;
	assign w30415 = w30450 ^ w30425;
	assign w30449 = w30415 ^ w30417;
	assign w30373 = w30450 ^ w30474;
	assign w30365 = w30412 ^ w30373;
	assign w30372 = w30402 ^ w30365;
	assign w30448 = w30369 ^ w30372;
	assign w30446 = w30415 ^ w30368;
	assign w30444 = w30365 ^ w30366;
	assign w30440 = w30446 & w30476;
	assign w30439 = w30449 & w30488;
	assign w30438 = w30459 & w30478;
	assign w30382 = w30438 ^ w30439;
	assign w30437 = w30447 & w30479;
	assign w30436 = w30444 & w30477;
	assign w30397 = w30436 ^ w30439;
	assign w30394 = ~w30397;
	assign w30393 = w30436 ^ w30437;
	assign w30435 = w30448 & w30480;
	assign w30431 = w30446 & w30491;
	assign w30413 = w30431 ^ w30435;
	assign w30398 = w30440 ^ w30431;
	assign w30391 = ~w30413;
	assign w30430 = w30449 & w30484;
	assign w30400 = w30438 ^ w30430;
	assign w30429 = w30459 & w30485;
	assign w30390 = w30391 ^ w30429;
	assign w30428 = w30447 & w30490;
	assign w30427 = w30444 & w30492;
	assign w30426 = w30448 & w30489;
	assign w30392 = w30437 ^ w30426;
	assign w30388 = ~w30392;
	assign w44644 = w30427 ^ w30428;
	assign w30409 = w30433 ^ w44644;
	assign w30410 = w30434 ^ w30409;
	assign w30414 = w30442 ^ w30410;
	assign w30383 = w30441 ^ w30414;
	assign w49860 = w30382 ^ w30383;
	assign w9074 = w9075 ^ w49860;
	assign w49735 = w9073 ^ w9074;
	assign w46849 = w49735 ^ w1073;
	assign w8890 = w49860 ^ w49850;
	assign w30419 = w30443 ^ w30414;
	assign w30494 = w30419 ^ w30393;
	assign w8972 = w30494 ^ w49853;
	assign w49862 = ~w30494;
	assign w9184 = w45348 ^ w49862;
	assign w9082 = w9192 ^ w9184;
	assign w9053 = w9184 ^ w9140;
	assign w49730 = w45610 ^ w9082;
	assign w49747 = w49858 ^ w9053;
	assign w46854 = w49730 ^ w1068;
	assign w46837 = w49747 ^ w1085;
	assign w8991 = w9184 ^ w45617;
	assign w9066 = w9190 ^ w30494;
	assign w49738 = w9066 ^ w9067;
	assign w46846 = w49738 ^ w1076;
	assign w30396 = w30400 ^ w44644;
	assign w30395 = w30391 ^ w30396;
	assign w30495 = w30394 ^ w30395;
	assign w44647 = w30439 ^ w30440;
	assign w49861 = w44647 ^ w30419;
	assign w8926 = w9141 ^ w49861;
	assign w9211 = w8926 ^ w8927;
	assign w49736 = w9211 ^ w9195;
	assign w46848 = w49736 ^ w1074;
	assign w16334 = w46848 ^ w46846;
	assign w9191 = w49857 ^ w49861;
	assign w9084 = w9086 ^ w9191;
	assign w9056 = w9192 ^ w9191;
	assign w49745 = w45347 ^ w9056;
	assign w46839 = w49745 ^ w1083;
	assign w9009 = w49861 ^ w12001;
	assign w30421 = w30436 ^ w44647;
	assign w30387 = w30432 ^ w30421;
	assign w30384 = ~w30387;
	assign w30381 = w30437 ^ w30421;
	assign w49863 = w30410 ^ w30381;
	assign w9147 = w49847 ^ w49863;
	assign w9132 = w9180 ^ w9147;
	assign w8889 = w9147 ^ w49845;
	assign w9226 = w8889 ^ w8890;
	assign w49720 = w9226 ^ w9191;
	assign w46864 = w49720 ^ w1058;
	assign w44648 = w30441 ^ w30443;
	assign w30399 = w44648 ^ w30396;
	assign w30496 = w30398 ^ w30399;
	assign w30386 = w30390 ^ w44648;
	assign w30389 = w30428 ^ w30386;
	assign w30493 = w30388 ^ w30389;
	assign w30385 = w30409 ^ w30386;
	assign w49859 = w30384 ^ w30385;
	assign w9182 = w49844 ^ w49859;
	assign w9044 = ~w9182;
	assign w9113 = w9044 ^ w45240;
	assign w49726 = w9113 ^ w9114;
	assign w9076 = w9182 ^ w9181;
	assign w49734 = w49848 ^ w9076;
	assign w46850 = w49734 ^ w1072;
	assign w16308 = w46849 ^ w46850;
	assign w16422 = w46850 ^ w46848;
	assign w17201 = w17223 & w17214;
	assign w44087 = w17201 ^ w17207;
	assign w17113 = w17145 ^ w44087;
	assign w17151 = w44087 ^ w17136;
	assign w17197 = w17159 ^ w17151;
	assign w44088 = w17201 ^ w17204;
	assign w17154 = w17202 ^ w44088;
	assign w17110 = w17205 ^ w17154;
	assign w17192 = w46995 ^ w17110;
	assign w17114 = w17140 ^ w44088;
	assign w17198 = w17114 ^ w17139;
	assign w17195 = w17196 ^ w17198;
	assign w17194 = w17197 & w17195;
	assign w17105 = w17194 ^ w17206;
	assign w17101 = w17105 ^ w17141;
	assign w17104 = w46989 ^ w17101;
	assign w17100 = w46991 ^ w17101;
	assign w17102 = w17194 ^ w17150;
	assign w17156 = w46991 ^ w17113;
	assign w17191 = w17196 ^ w17156;
	assign w17190 = w17191 & w17192;
	assign w17189 = w17190 ^ w17198;
	assign w17166 = w17189 & w17221;
	assign w17108 = w17190 ^ w17207;
	assign w17103 = w17108 ^ w17204;
	assign w17181 = w17103 ^ w17104;
	assign w17193 = w17194 ^ w17156;
	assign w17109 = w17190 ^ w17154;
	assign w17162 = w17181 & w17224;
	assign w17163 = w17193 & w17219;
	assign w17175 = w17189 & w46996;
	assign w17172 = w17193 & w17212;
	assign w17171 = w17181 & w17213;
	assign w17188 = w17196 ^ w17190;
	assign w17187 = w17198 & w17188;
	assign w17185 = w17187 ^ w17195;
	assign w17184 = w17193 & w17185;
	assign w17107 = w17184 ^ w17208;
	assign w17149 = w17184 ^ w17159;
	assign w17183 = w17149 ^ w17151;
	assign w17180 = w17149 ^ w17102;
	assign w17174 = w17180 & w17210;
	assign w17173 = w17183 & w17222;
	assign w17116 = w17172 ^ w17173;
	assign w17165 = w17180 & w17225;
	assign w17132 = w17174 ^ w17165;
	assign w17164 = w17183 & w17218;
	assign w17134 = w17172 ^ w17164;
	assign w44089 = w17173 ^ w17174;
	assign w44091 = w17187 ^ w17205;
	assign w17179 = w44091 ^ w17157;
	assign w17177 = w17179 & w17216;
	assign w44090 = w17175 ^ w17177;
	assign w17168 = w17179 & w17220;
	assign w17146 = w46995 ^ w44091;
	assign w17186 = w17146 ^ w17109;
	assign w17176 = w17186 & w17215;
	assign w17099 = w17146 ^ w17107;
	assign w17106 = w17136 ^ w17099;
	assign w17182 = w17103 ^ w17106;
	assign w17178 = w17099 ^ w17100;
	assign w17170 = w17178 & w17211;
	assign w17155 = w17170 ^ w44089;
	assign w17131 = w17170 ^ w17173;
	assign w17128 = ~w17131;
	assign w17127 = w17170 ^ w17171;
	assign w17121 = w17166 ^ w17155;
	assign w17118 = ~w17121;
	assign w17169 = w17182 & w17214;
	assign w17147 = w17165 ^ w17169;
	assign w17125 = ~w17147;
	assign w17124 = w17125 ^ w17163;
	assign w17120 = w17124 ^ w44090;
	assign w17123 = w17162 ^ w17120;
	assign w17161 = w17178 & w17226;
	assign w43546 = w17161 ^ w17162;
	assign w17130 = w17134 ^ w43546;
	assign w17129 = w17125 ^ w17130;
	assign w17229 = w17128 ^ w17129;
	assign w17133 = w44090 ^ w17130;
	assign w17230 = w17132 ^ w17133;
	assign w17167 = w17186 & w17217;
	assign w17143 = w17167 ^ w43546;
	assign w17144 = w17168 ^ w17143;
	assign w17119 = w17143 ^ w17120;
	assign w17148 = w17176 ^ w17144;
	assign w17117 = w17175 ^ w17148;
	assign w49901 = w17116 ^ w17117;
	assign w17153 = w17177 ^ w17148;
	assign w49902 = w44089 ^ w17153;
	assign w17228 = w17153 ^ w17127;
	assign w9159 = w49901 ^ w49914;
	assign w8939 = ~w49902;
	assign w9093 = w9229 ^ w49901;
	assign w9128 = w49915 ^ w8939;
	assign w49903 = ~w17228;
	assign w9130 = w9159 ^ w9150;
	assign w49900 = w17118 ^ w17119;
	assign w17115 = w17171 ^ w17155;
	assign w49904 = w17144 ^ w17115;
	assign w9145 = w49904 ^ w49916;
	assign w8944 = w9183 ^ w9145;
	assign w8901 = w9145 ^ w49900;
	assign w9221 = w8901 ^ w8902;
	assign w9194 = w49856 ^ w49860;
	assign w9059 = w9195 ^ w9194;
	assign w49727 = w9209 ^ w9194;
	assign w9057 = ~w9059;
	assign w46857 = w49727 ^ w1065;
	assign w9041 = w9194 ^ w9044;
	assign w9139 = w49858 ^ w49863;
	assign w9063 = w9180 ^ w9139;
	assign w49740 = w45612 ^ w9063;
	assign w46844 = w49740 ^ w1078;
	assign w9081 = w9190 ^ w9139;
	assign w49731 = w49847 ^ w9081;
	assign w46853 = w49731 ^ w1069;
	assign w9043 = ~w9147;
	assign w9042 = w9043 ^ w49849;
	assign w49719 = w9041 ^ w9042;
	assign w17160 = w17182 & w17223;
	assign w17126 = w17171 ^ w17160;
	assign w17122 = ~w17126;
	assign w17227 = w17122 ^ w17123;
	assign w46865 = w49719 ^ w1057;
	assign w46858 = w49726 ^ w1064;
	assign w11752 = w46857 ^ w46858;
	assign w11863 = w46853 ^ w46858;
	assign w45362 = ~w17230;
	assign w8899 = w9145 ^ w45362;
	assign w45368 = ~w17227;
	assign w9112 = w17228 ^ w45368;
	assign w9168 = w45368 ^ w45690;
	assign w9102 = w9168 ^ w49911;
	assign w9126 = w9168 ^ w9156;
	assign w45369 = ~w17229;
	assign w8942 = w9151 ^ w45369;
	assign w23970 = w46839 ^ w46837;
	assign w45699 = ~w30493;
	assign w9068 = w9192 ^ w45699;
	assign w49737 = w9068 ^ w9069;
	assign w46847 = w49737 ^ w1075;
	assign w16293 = w16334 ^ w46847;
	assign w9187 = w45347 ^ w45699;
	assign w9083 = w9195 ^ w9187;
	assign w49729 = w45617 ^ w9083;
	assign w9054 = w9190 ^ w9187;
	assign w46855 = w49729 ^ w1067;
	assign w11776 = w46855 ^ w46853;
	assign w9010 = w9187 ^ w49846;
	assign w9008 = ~w9010;
	assign w49721 = w9008 ^ w9009;
	assign w46863 = w49721 ^ w1059;
	assign w8992 = w45699 ^ w12002;
	assign w8990 = w8991 ^ w8992;
	assign w49722 = ~w8990;
	assign w46862 = w49722 ^ w1060;
	assign w27054 = w46864 ^ w46862;
	assign w27013 = w27054 ^ w46863;
	assign w49746 = w45348 ^ w9054;
	assign w46838 = w49746 ^ w1084;
	assign w23976 = w46844 ^ w46838;
	assign w24053 = w23970 ^ w23976;
	assign w24056 = w46839 ^ w23976;
	assign w45700 = ~w30495;
	assign w9061 = w45700 ^ w16559;
	assign w49742 = w9060 ^ w9061;
	assign w46842 = w49742 ^ w1080;
	assign w24057 = w46837 ^ w46842;
	assign w9202 = w45611 ^ w45700;
	assign w9078 = w9202 ^ w9180;
	assign w9055 = w9202 ^ w9179;
	assign w9077 = w9078 ^ w9079;
	assign w49733 = ~w9077;
	assign w46851 = w49733 ^ w1071;
	assign w16348 = w46851 ^ w46850;
	assign w49718 = w49859 ^ w9055;
	assign w46866 = w49718 ^ w1056;
	assign w27142 = w46866 ^ w46864;
	assign w27028 = w46865 ^ w46866;
	assign w16331 = w46851 ^ w46849;
	assign w16333 = w46850 ^ w16331;
	assign w16409 = w46846 ^ w16333;
	assign w16406 = w46847 ^ w16333;
	assign w45701 = ~w30496;
	assign w8932 = w9139 ^ w45701;
	assign w9203 = w45612 ^ w45701;
	assign w9080 = w9203 ^ w9141;
	assign w49732 = w45241 ^ w9080;
	assign w46852 = w49732 ^ w1070;
	assign w16417 = w46852 ^ w16293;
	assign w16403 = w46852 & w16417;
	assign w9071 = w9203 ^ w9181;
	assign w49716 = w45701 ^ w9132;
	assign w46868 = w49716 ^ w1054;
	assign w27058 = w46868 ^ w46862;
	assign w27138 = w46863 ^ w27058;
	assign w27137 = w46868 ^ w27013;
	assign w27123 = w46868 & w27137;
	assign w8955 = w9203 ^ w9140;
	assign w49724 = w45349 ^ w8955;
	assign w46860 = w49724 ^ w1062;
	assign w11782 = w46860 ^ w46854;
	assign w11862 = w46855 ^ w11782;
	assign w11859 = w11776 ^ w11782;
	assign w9208 = w8932 ^ w8933;
	assign w49741 = w9208 ^ w9181;
	assign w46843 = w49741 ^ w1079;
	assign w24059 = w46837 ^ w46843;
	assign w16338 = w46852 ^ w46846;
	assign w16418 = w46847 ^ w16338;
	assign w16414 = w46851 ^ w16418;
	assign w16401 = w16418 & w16414;
	assign w23986 = w46843 ^ w46842;
	assign w24051 = w23986 ^ w24053;
	assign w24052 = w46843 ^ w24056;
	assign w24039 = w24056 & w24052;
	assign w16408 = w16338 ^ w16333;
	assign w9072 = w9043 ^ w45700;
	assign w9070 = w9071 ^ w9072;
	assign w49717 = ~w9070;
	assign w46867 = w49717 ^ w1055;
	assign w27051 = w46867 ^ w46865;
	assign w27053 = w46866 ^ w27051;
	assign w27068 = w46867 ^ w46866;
	assign w27134 = w46867 ^ w27138;
	assign w27121 = w27138 & w27134;
	assign w27129 = w46862 ^ w27053;
	assign w27126 = w46863 ^ w27053;
	assign w27128 = w27058 ^ w27053;
	assign w45938 = ~w8793;
	assign w8691 = w45938 ^ w49664;
	assign w49558 = w8690 ^ w8691;
	assign w8688 = w45938 ^ w49665;
	assign w49559 = w8687 ^ w8688;
	assign w8695 = w45938 ^ w45615;
	assign w46953 = w49558 ^ w906;
	assign w12020 = w46953 ^ w46954;
	assign w46952 = w49559 ^ w907;
	assign w12134 = w46954 ^ w46952;
	assign w12132 = w46952 ^ w46949;
	assign w12119 = w12044 ^ w12134;
	assign w12110 = w12134 & w12119;
	assign w12046 = w46952 ^ w46950;
	assign w12006 = w12046 ^ w12044;
	assign w12005 = w12046 ^ w46951;
	assign w12129 = w46956 ^ w12005;
	assign w12115 = w46956 & w12129;
	assign w8693 = w8694 ^ w8695;
	assign w49556 = ~w8693;
	assign w46955 = w49556 ^ w904;
	assign w12060 = w46955 ^ w46954;
	assign w12128 = w12132 ^ w12060;
	assign w12125 = w12060 ^ w12127;
	assign w12043 = w46955 ^ w46953;
	assign w12122 = w12043 ^ w12006;
	assign w12109 = w12131 & w12122;
	assign w12045 = w46954 ^ w12043;
	assign w12118 = w46951 ^ w12045;
	assign w12120 = w12050 ^ w12045;
	assign w12112 = w12127 & w12120;
	assign w12121 = w46950 ^ w12045;
	assign w12111 = w12132 & w12121;
	assign w12047 = w12111 ^ w12045;
	assign w12133 = w46949 ^ w46955;
	assign w12114 = w12133 & w12118;
	assign w12048 = w12114 ^ w12044;
	assign w12126 = w46955 ^ w12130;
	assign w12113 = w12130 & w12126;
	assign w12124 = w12043 ^ w12132;
	assign w12117 = w12124 & w12128;
	assign w12049 = w12117 ^ w12046;
	assign w12053 = w12049 ^ w12047;
	assign w12058 = w46949 ^ w12053;
	assign w12123 = w46956 ^ w12124;
	assign w43875 = w12109 ^ w12115;
	assign w12059 = w43875 ^ w12044;
	assign w12021 = w12053 ^ w43875;
	assign w12064 = w46951 ^ w12021;
	assign w43876 = w12109 ^ w12112;
	assign w12062 = w12110 ^ w43876;
	assign w12018 = w12113 ^ w12062;
	assign w12100 = w46955 ^ w12018;
	assign w12022 = w12048 ^ w43876;
	assign w12106 = w12022 ^ w12047;
	assign w12019 = w12110 ^ w12111;
	assign w12066 = w12019 ^ w12020;
	assign w12065 = w12066 ^ w12048;
	assign w12107 = w12113 ^ w12065;
	assign w12116 = w12125 & w12123;
	assign w12067 = w12110 ^ w12116;
	assign w12105 = w12067 ^ w12059;
	assign w12108 = w12067 ^ w12058;
	assign w12104 = w12108 & w12107;
	assign w12103 = w12104 ^ w12106;
	assign w12102 = w12105 & w12103;
	assign w12010 = w12102 ^ w12058;
	assign w12101 = w12102 ^ w12064;
	assign w12071 = w12101 & w12127;
	assign w12099 = w12104 ^ w12064;
	assign w12098 = w12099 & w12100;
	assign w12016 = w12098 ^ w12115;
	assign w12011 = w12016 ^ w12112;
	assign w12017 = w12098 ^ w12062;
	assign w12096 = w12104 ^ w12098;
	assign w12095 = w12106 & w12096;
	assign w12093 = w12095 ^ w12103;
	assign w12092 = w12101 & w12093;
	assign w12057 = w12092 ^ w12067;
	assign w12088 = w12057 ^ w12010;
	assign w12091 = w12057 ^ w12059;
	assign w12081 = w12091 & w12130;
	assign w12072 = w12091 & w12126;
	assign w12013 = w12102 ^ w12114;
	assign w12009 = w12013 ^ w12049;
	assign w12008 = w46951 ^ w12009;
	assign w12012 = w46949 ^ w12009;
	assign w12089 = w12011 ^ w12012;
	assign w12070 = w12089 & w12132;
	assign w43879 = w12095 ^ w12113;
	assign w12054 = w46955 ^ w43879;
	assign w12094 = w12054 ^ w12017;
	assign w12084 = w12094 & w12123;
	assign w12075 = w12094 & w12125;
	assign w12087 = w43879 ^ w12065;
	assign w12076 = w12087 & w12128;
	assign w12085 = w12087 & w12124;
	assign w12015 = w12092 ^ w12116;
	assign w12007 = w12054 ^ w12015;
	assign w12014 = w12044 ^ w12007;
	assign w12086 = w12007 ^ w12008;
	assign w12090 = w12011 ^ w12014;
	assign w12077 = w12090 & w12122;
	assign w12068 = w12090 & w12131;
	assign w12097 = w12098 ^ w12106;
	assign w12083 = w12097 & w46956;
	assign w12074 = w12097 & w12129;
	assign w43878 = w12083 ^ w12085;
	assign w12082 = w12088 & w12118;
	assign w43877 = w12081 ^ w12082;
	assign w12069 = w12086 & w12134;
	assign w43530 = w12069 ^ w12070;
	assign w12051 = w12075 ^ w43530;
	assign w12052 = w12076 ^ w12051;
	assign w12056 = w12084 ^ w12052;
	assign w12061 = w12085 ^ w12056;
	assign w49907 = w43877 ^ w12061;
	assign w9199 = w49902 ^ w49907;
	assign w49840 = w9205 ^ w9199;
	assign w9115 = w9199 ^ w9168;
	assign w49825 = w45613 ^ w9115;
	assign w12025 = w12083 ^ w12056;
	assign w46759 = w49825 ^ w972;
	assign w46744 = w49840 ^ w986;
	assign w9131 = w9145 ^ w49907;
	assign w49816 = w9130 ^ w9131;
	assign w46768 = w49816 ^ w963;
	assign w12080 = w12101 & w12120;
	assign w12042 = w12080 ^ w12072;
	assign w12024 = w12080 ^ w12081;
	assign w12038 = w12042 ^ w43530;
	assign w12041 = w43878 ^ w12038;
	assign w49906 = w12024 ^ w12025;
	assign w9153 = w49906 ^ w49910;
	assign w49815 = w9221 ^ w9153;
	assign w9092 = w9153 ^ w9151;
	assign w9104 = w9199 ^ w9153;
	assign w9091 = w9092 ^ w9093;
	assign w49839 = ~w9091;
	assign w46769 = w49815 ^ w962;
	assign w8938 = w49906 ^ w8939;
	assign w46745 = w49839 ^ w45170;
	assign w12079 = w12089 & w12121;
	assign w12034 = w12079 ^ w12068;
	assign w12030 = ~w12034;
	assign w12078 = w12086 & w12119;
	assign w12063 = w12078 ^ w43877;
	assign w12039 = w12078 ^ w12081;
	assign w12036 = ~w12039;
	assign w12023 = w12079 ^ w12063;
	assign w49908 = w12052 ^ w12023;
	assign w9148 = w49908 ^ w49912;
	assign w9134 = w49904 ^ w49908;
	assign w9099 = w9134 ^ w49916;
	assign w9123 = w9183 ^ w9134;
	assign w9087 = w9156 ^ w9134;
	assign w9125 = w49908 ^ w17228;
	assign w49819 = w9124 ^ w9125;
	assign w49820 = w45362 ^ w9123;
	assign w49843 = w49912 ^ w9087;
	assign w46741 = w49843 ^ w989;
	assign w23924 = w46744 ^ w46741;
	assign w46764 = w49820 ^ w967;
	assign w46765 = w49819 ^ w966;
	assign w26872 = w46768 ^ w46765;
	assign w12035 = w12078 ^ w12079;
	assign w12136 = w12061 ^ w12035;
	assign w8887 = w9148 ^ w49909;
	assign w8885 = w9148 ^ w45692;
	assign w9105 = w9148 ^ w49915;
	assign w49832 = w9104 ^ w9105;
	assign w46752 = w49832 ^ w979;
	assign w12029 = w12074 ^ w12063;
	assign w12026 = ~w12029;
	assign w45245 = ~w12136;
	assign w9100 = w45606 ^ w45245;
	assign w9198 = w49903 ^ w45245;
	assign w9088 = w9198 ^ w45690;
	assign w49842 = w9088 ^ w9089;
	assign w49818 = w45245 ^ w9126;
	assign w9109 = w9198 ^ w9133;
	assign w49827 = w49904 ^ w9109;
	assign w49835 = w9099 ^ w9100;
	assign w46757 = w49827 ^ w974;
	assign w11508 = w46759 ^ w46757;
	assign w46749 = w49835 ^ w982;
	assign w46766 = w49818 ^ w965;
	assign w46742 = w49842 ^ w988;
	assign w23838 = w46744 ^ w46742;
	assign w15884 = w46752 ^ w46749;
	assign w26786 = w46768 ^ w46766;
	assign w12073 = w12088 & w12133;
	assign w12055 = w12073 ^ w12077;
	assign w12040 = w12082 ^ w12073;
	assign w12138 = w12040 ^ w12041;
	assign w12033 = ~w12055;
	assign w12037 = w12033 ^ w12038;
	assign w12032 = w12033 ^ w12071;
	assign w12028 = w12032 ^ w43878;
	assign w12031 = w12070 ^ w12028;
	assign w12135 = w12030 ^ w12031;
	assign w12027 = w12051 ^ w12028;
	assign w49905 = w12026 ^ w12027;
	assign w9173 = w49900 ^ w49905;
	assign w9094 = w9173 ^ w9163;
	assign w9118 = w9173 ^ w9159;
	assign w9116 = ~w9118;
	assign w49838 = w49909 ^ w9094;
	assign w9106 = w9173 ^ w49913;
	assign w46746 = w49838 ^ w985;
	assign w23812 = w46745 ^ w46746;
	assign w23923 = w46741 ^ w46746;
	assign w8888 = w49906 ^ w49905;
	assign w9227 = w8887 ^ w8888;
	assign w49831 = w9227 ^ w9159;
	assign w46753 = w49831 ^ w978;
	assign w8943 = w45692 ^ w49905;
	assign w49814 = w8942 ^ w8943;
	assign w46770 = w49814 ^ w961;
	assign w26760 = w46769 ^ w46770;
	assign w26871 = w46765 ^ w46770;
	assign w45239 = ~w12138;
	assign w9196 = w45362 ^ w45239;
	assign w9121 = w9196 ^ w9163;
	assign w9098 = w9196 ^ w9133;
	assign w49836 = w45608 ^ w9098;
	assign w9108 = w9196 ^ w9148;
	assign w49828 = w45693 ^ w9108;
	assign w46756 = w49828 ^ w975;
	assign w8886 = w45608 ^ w45239;
	assign w9228 = w8885 ^ w8886;
	assign w46748 = w49836 ^ w983;
	assign w23842 = w46748 ^ w46742;
	assign w49812 = w45239 ^ w8944;
	assign w46772 = w49812 ^ w959;
	assign w26790 = w46772 ^ w46766;
	assign w45244 = ~w12135;
	assign w9158 = w45244 ^ w45613;
	assign w9111 = w9156 ^ w45244;
	assign w9101 = w9198 ^ w9158;
	assign w49834 = w45691 ^ w9101;
	assign w9090 = w9158 ^ w9150;
	assign w9103 = w45244 ^ w49907;
	assign w49833 = w9102 ^ w9103;
	assign w9110 = w9111 ^ w9112;
	assign w49826 = ~w9110;
	assign w46758 = w49826 ^ w973;
	assign w46751 = w49833 ^ w980;
	assign w15796 = w46751 ^ w46749;
	assign w9129 = ~w9158;
	assign w11514 = w46764 ^ w46758;
	assign w11591 = w11508 ^ w11514;
	assign w46750 = w49834 ^ w981;
	assign w15802 = w46756 ^ w46750;
	assign w15798 = w46752 ^ w46750;
	assign w15879 = w15796 ^ w15802;
	assign w15882 = w46751 ^ w15802;
	assign w15757 = w15798 ^ w46751;
	assign w15881 = w46756 ^ w15757;
	assign w11594 = w46759 ^ w11514;
	assign w49841 = w45368 ^ w9090;
	assign w46743 = w49841 ^ w987;
	assign w23836 = w46743 ^ w46741;
	assign w23798 = w23838 ^ w23836;
	assign w23922 = w46743 ^ w23842;
	assign w23919 = w23836 ^ w23842;
	assign w23797 = w23838 ^ w46743;
	assign w23921 = w46748 ^ w23797;
	assign w23907 = w46748 & w23921;
	assign w9127 = w9129 ^ w45690;
	assign w49817 = w9127 ^ w9128;
	assign w46767 = w49817 ^ w964;
	assign w26784 = w46767 ^ w46765;
	assign w26867 = w26784 ^ w26790;
	assign w26746 = w26786 ^ w26784;
	assign w26745 = w26786 ^ w46767;
	assign w26869 = w46772 ^ w26745;
	assign w26855 = w46772 & w26869;
	assign w23926 = w46746 ^ w46744;
	assign w23911 = w23836 ^ w23926;
	assign w23902 = w23926 & w23911;
	assign w12137 = w12036 ^ w12037;
	assign w45238 = ~w12137;
	assign w9107 = w45607 ^ w45238;
	assign w49830 = w9106 ^ w9107;
	assign w46754 = w49830 ^ w977;
	assign w15886 = w46754 ^ w46752;
	assign w15883 = w46749 ^ w46754;
	assign w15772 = w46753 ^ w46754;
	assign w15871 = w15796 ^ w15886;
	assign w15862 = w15886 & w15871;
	assign w9188 = w45369 ^ w45238;
	assign w9119 = w9188 ^ w9151;
	assign w49829 = w9228 ^ w9188;
	assign w9097 = ~w9188;
	assign w49822 = w49900 ^ w9119;
	assign w9095 = w9097 ^ w9183;
	assign w49837 = w9095 ^ w9096;
	assign w46762 = w49822 ^ w969;
	assign w11595 = w46757 ^ w46762;
	assign w46747 = w49837 ^ w984;
	assign w46755 = w49829 ^ w976;
	assign w15878 = w46755 ^ w15882;
	assign w15885 = w46749 ^ w46755;
	assign w15795 = w46755 ^ w46753;
	assign w15876 = w15795 ^ w15884;
	assign w15875 = w46756 ^ w15876;
	assign w15865 = w15882 & w15878;
	assign w15812 = w46755 ^ w46754;
	assign w15880 = w15884 ^ w15812;
	assign w15869 = w15876 & w15880;
	assign w15877 = w15812 ^ w15879;
	assign w15868 = w15877 & w15875;
	assign w23918 = w46747 ^ w23922;
	assign w23905 = w23922 & w23918;
	assign w15797 = w46754 ^ w15795;
	assign w15873 = w46750 ^ w15797;
	assign w15870 = w46751 ^ w15797;
	assign w15866 = w15885 & w15870;
	assign w15863 = w15884 & w15873;
	assign w15771 = w15862 ^ w15863;
	assign w15818 = w15771 ^ w15772;
	assign w15872 = w15802 ^ w15797;
	assign w15864 = w15879 & w15872;
	assign w15800 = w15866 ^ w15796;
	assign w15799 = w15863 ^ w15797;
	assign w15801 = w15869 ^ w15798;
	assign w15805 = w15801 ^ w15799;
	assign w15810 = w46749 ^ w15805;
	assign w15819 = w15862 ^ w15868;
	assign w15860 = w15819 ^ w15810;
	assign w8900 = w45693 ^ w45238;
	assign w23925 = w46741 ^ w46747;
	assign w15817 = w15818 ^ w15800;
	assign w15859 = w15865 ^ w15817;
	assign w15856 = w15860 & w15859;
	assign w9222 = w8899 ^ w8900;
	assign w49813 = w9222 ^ w9163;
	assign w46771 = w49813 ^ w960;
	assign w26873 = w46765 ^ w46771;
	assign w26783 = w46771 ^ w46769;
	assign w26785 = w46770 ^ w26783;
	assign w26858 = w46767 ^ w26785;
	assign w26854 = w26873 & w26858;
	assign w26860 = w26790 ^ w26785;
	assign w26852 = w26867 & w26860;
	assign w26862 = w26783 ^ w26746;
	assign w26849 = w26871 & w26862;
	assign w26864 = w26783 ^ w26872;
	assign w26863 = w46772 ^ w26864;
	assign w26861 = w46766 ^ w26785;
	assign w26851 = w26872 & w26861;
	assign w26787 = w26851 ^ w26785;
	assign w44493 = w26849 ^ w26855;
	assign w26799 = w44493 ^ w26784;
	assign w26788 = w26854 ^ w26784;
	assign w44490 = w26849 ^ w26852;
	assign w26762 = w26788 ^ w44490;
	assign w26846 = w26762 ^ w26787;
	assign w26800 = w46771 ^ w46770;
	assign w26868 = w26872 ^ w26800;
	assign w26857 = w26864 & w26868;
	assign w26789 = w26857 ^ w26786;
	assign w26793 = w26789 ^ w26787;
	assign w26798 = w46765 ^ w26793;
	assign w26761 = w26793 ^ w44493;
	assign w26804 = w46767 ^ w26761;
	assign w26865 = w26800 ^ w26867;
	assign w26856 = w26865 & w26863;
	assign w23835 = w46747 ^ w46745;
	assign w23837 = w46746 ^ w23835;
	assign w23912 = w23842 ^ w23837;
	assign w23904 = w23919 & w23912;
	assign w23910 = w46743 ^ w23837;
	assign w23914 = w23835 ^ w23798;
	assign w23901 = w23923 & w23914;
	assign w23916 = w23835 ^ w23924;
	assign w23915 = w46748 ^ w23916;
	assign w44368 = w23901 ^ w23907;
	assign w23851 = w44368 ^ w23836;
	assign w44369 = w23901 ^ w23904;
	assign w23854 = w23902 ^ w44369;
	assign w23810 = w23905 ^ w23854;
	assign w23892 = w46747 ^ w23810;
	assign w23913 = w46742 ^ w23837;
	assign w23903 = w23924 & w23913;
	assign w23839 = w23903 ^ w23837;
	assign w23811 = w23902 ^ w23903;
	assign w23858 = w23811 ^ w23812;
	assign w23906 = w23925 & w23910;
	assign w23840 = w23906 ^ w23836;
	assign w23814 = w23840 ^ w44369;
	assign w23898 = w23814 ^ w23839;
	assign w23857 = w23858 ^ w23840;
	assign w23899 = w23905 ^ w23857;
	assign w23852 = w46747 ^ w46746;
	assign w23917 = w23852 ^ w23919;
	assign w23908 = w23917 & w23915;
	assign w23920 = w23924 ^ w23852;
	assign w23859 = w23902 ^ w23908;
	assign w23897 = w23859 ^ w23851;
	assign w23909 = w23916 & w23920;
	assign w23841 = w23909 ^ w23838;
	assign w23845 = w23841 ^ w23839;
	assign w23813 = w23845 ^ w44368;
	assign w23856 = w46743 ^ w23813;
	assign w23850 = w46741 ^ w23845;
	assign w23900 = w23859 ^ w23850;
	assign w23896 = w23900 & w23899;
	assign w23891 = w23896 ^ w23856;
	assign w23890 = w23891 & w23892;
	assign w23889 = w23890 ^ w23898;
	assign w23808 = w23890 ^ w23907;
	assign w23803 = w23808 ^ w23904;
	assign w23875 = w23889 & w46748;
	assign w23888 = w23896 ^ w23890;
	assign w23887 = w23898 & w23888;
	assign w23895 = w23896 ^ w23898;
	assign w23885 = w23887 ^ w23895;
	assign w23894 = w23897 & w23895;
	assign w23802 = w23894 ^ w23850;
	assign w23805 = w23894 ^ w23906;
	assign w23801 = w23805 ^ w23841;
	assign w23800 = w46743 ^ w23801;
	assign w23893 = w23894 ^ w23856;
	assign w23863 = w23893 & w23919;
	assign w23872 = w23893 & w23912;
	assign w23884 = w23893 & w23885;
	assign w23807 = w23884 ^ w23908;
	assign w23849 = w23884 ^ w23859;
	assign w23880 = w23849 ^ w23802;
	assign w23874 = w23880 & w23910;
	assign w23883 = w23849 ^ w23851;
	assign w23864 = w23883 & w23918;
	assign w23834 = w23872 ^ w23864;
	assign w23873 = w23883 & w23922;
	assign w23816 = w23872 ^ w23873;
	assign w44371 = w23873 ^ w23874;
	assign w44373 = w23887 ^ w23905;
	assign w23879 = w44373 ^ w23857;
	assign w23877 = w23879 & w23916;
	assign w23868 = w23879 & w23920;
	assign w44372 = w23875 ^ w23877;
	assign w23804 = w46741 ^ w23801;
	assign w23881 = w23803 ^ w23804;
	assign w23862 = w23881 & w23924;
	assign w23871 = w23881 & w23913;
	assign w23866 = w23889 & w23921;
	assign w23846 = w46747 ^ w44373;
	assign w23799 = w23846 ^ w23807;
	assign w23806 = w23836 ^ w23799;
	assign w23882 = w23803 ^ w23806;
	assign w23860 = w23882 & w23923;
	assign w23869 = w23882 & w23914;
	assign w23826 = w23871 ^ w23860;
	assign w23822 = ~w23826;
	assign w23878 = w23799 ^ w23800;
	assign w23870 = w23878 & w23911;
	assign w23855 = w23870 ^ w44371;
	assign w23821 = w23866 ^ w23855;
	assign w23815 = w23871 ^ w23855;
	assign w23818 = ~w23821;
	assign w23827 = w23870 ^ w23871;
	assign w23861 = w23878 & w23926;
	assign w23831 = w23870 ^ w23873;
	assign w23828 = ~w23831;
	assign w44370 = w23861 ^ w23862;
	assign w23830 = w23834 ^ w44370;
	assign w23833 = w44372 ^ w23830;
	assign w23865 = w23880 & w23925;
	assign w23832 = w23874 ^ w23865;
	assign w23930 = w23832 ^ w23833;
	assign w23847 = w23865 ^ w23869;
	assign w23825 = ~w23847;
	assign w23824 = w23825 ^ w23863;
	assign w23820 = w23824 ^ w44372;
	assign w23823 = w23862 ^ w23820;
	assign w23809 = w23890 ^ w23854;
	assign w45516 = ~w23930;
	assign w9528 = w45333 ^ w45516;
	assign w26874 = w46770 ^ w46768;
	assign w26859 = w26784 ^ w26874;
	assign w26850 = w26874 & w26859;
	assign w26802 = w26850 ^ w44490;
	assign w26759 = w26850 ^ w26851;
	assign w26806 = w26759 ^ w26760;
	assign w26805 = w26806 ^ w26788;
	assign w26807 = w26850 ^ w26856;
	assign w26848 = w26807 ^ w26798;
	assign w26845 = w26807 ^ w26799;
	assign w26870 = w46767 ^ w26790;
	assign w26866 = w46771 ^ w26870;
	assign w26853 = w26870 & w26866;
	assign w26847 = w26853 ^ w26805;
	assign w26758 = w26853 ^ w26802;
	assign w26840 = w46771 ^ w26758;
	assign w26844 = w26848 & w26847;
	assign w26839 = w26844 ^ w26804;
	assign w26838 = w26839 & w26840;
	assign w26757 = w26838 ^ w26802;
	assign w26756 = w26838 ^ w26855;
	assign w26836 = w26844 ^ w26838;
	assign w26751 = w26756 ^ w26852;
	assign w26835 = w26846 & w26836;
	assign w44492 = w26835 ^ w26853;
	assign w26827 = w44492 ^ w26805;
	assign w26816 = w26827 & w26868;
	assign w26825 = w26827 & w26864;
	assign w26794 = w46771 ^ w44492;
	assign w26834 = w26794 ^ w26757;
	assign w26824 = w26834 & w26863;
	assign w26815 = w26834 & w26865;
	assign w26837 = w26838 ^ w26846;
	assign w26823 = w26837 & w46772;
	assign w26814 = w26837 & w26869;
	assign w44495 = w26823 ^ w26825;
	assign w26843 = w26844 ^ w26846;
	assign w26833 = w26835 ^ w26843;
	assign w26842 = w26845 & w26843;
	assign w26841 = w26842 ^ w26804;
	assign w26832 = w26841 & w26833;
	assign w26755 = w26832 ^ w26856;
	assign w26747 = w26794 ^ w26755;
	assign w26754 = w26784 ^ w26747;
	assign w26830 = w26751 ^ w26754;
	assign w26820 = w26841 & w26860;
	assign w26797 = w26832 ^ w26807;
	assign w26753 = w26842 ^ w26854;
	assign w26749 = w26753 ^ w26789;
	assign w26748 = w46767 ^ w26749;
	assign w26826 = w26747 ^ w26748;
	assign w26817 = w26830 & w26862;
	assign w26752 = w46765 ^ w26749;
	assign w26829 = w26751 ^ w26752;
	assign w26810 = w26829 & w26872;
	assign w26819 = w26829 & w26861;
	assign w26831 = w26797 ^ w26799;
	assign w26750 = w26842 ^ w26798;
	assign w26828 = w26797 ^ w26750;
	assign w26822 = w26828 & w26858;
	assign w26809 = w26826 & w26874;
	assign w26821 = w26831 & w26870;
	assign w26764 = w26820 ^ w26821;
	assign w26818 = w26826 & w26859;
	assign w26779 = w26818 ^ w26821;
	assign w26776 = ~w26779;
	assign w26775 = w26818 ^ w26819;
	assign w44491 = w26809 ^ w26810;
	assign w26791 = w26815 ^ w44491;
	assign w26792 = w26816 ^ w26791;
	assign w44494 = w26821 ^ w26822;
	assign w26796 = w26824 ^ w26792;
	assign w26765 = w26823 ^ w26796;
	assign w50083 = w26764 ^ w26765;
	assign w26813 = w26828 & w26873;
	assign w26780 = w26822 ^ w26813;
	assign w26795 = w26813 ^ w26817;
	assign w26773 = ~w26795;
	assign w26812 = w26831 & w26866;
	assign w26782 = w26820 ^ w26812;
	assign w26778 = w26782 ^ w44491;
	assign w26781 = w44495 ^ w26778;
	assign w26777 = w26773 ^ w26778;
	assign w26878 = w26780 ^ w26781;
	assign w26877 = w26776 ^ w26777;
	assign w26811 = w26841 & w26867;
	assign w26772 = w26773 ^ w26811;
	assign w26768 = w26772 ^ w44495;
	assign w26771 = w26810 ^ w26768;
	assign w26767 = w26791 ^ w26768;
	assign w45594 = ~w26877;
	assign w45595 = ~w26878;
	assign w26801 = w26825 ^ w26796;
	assign w50084 = w44494 ^ w26801;
	assign w26876 = w26801 ^ w26775;
	assign w45601 = ~w26876;
	assign w23927 = w23822 ^ w23823;
	assign w45521 = ~w23927;
	assign w15758 = w15798 ^ w15796;
	assign w15874 = w15795 ^ w15758;
	assign w15861 = w15883 & w15874;
	assign w44031 = w15861 ^ w15864;
	assign w15814 = w15862 ^ w44031;
	assign w15770 = w15865 ^ w15814;
	assign w15852 = w46755 ^ w15770;
	assign w15774 = w15800 ^ w44031;
	assign w15858 = w15774 ^ w15799;
	assign w15855 = w15856 ^ w15858;
	assign w23886 = w23846 ^ w23809;
	assign w23867 = w23886 & w23917;
	assign w23843 = w23867 ^ w44370;
	assign w23819 = w23843 ^ w23820;
	assign w23876 = w23886 & w23915;
	assign w23844 = w23868 ^ w23843;
	assign w50117 = w23844 ^ w23815;
	assign w23848 = w23876 ^ w23844;
	assign w23817 = w23875 ^ w23848;
	assign w50115 = w23816 ^ w23817;
	assign w23853 = w23877 ^ w23848;
	assign w50116 = w44371 ^ w23853;
	assign w9495 = w50112 ^ w50116;
	assign w23928 = w23853 ^ w23827;
	assign w9478 = w50113 ^ w50117;
	assign w9285 = w9478 ^ w50115;
	assign w9550 = w9285 ^ w9286;
	assign w50114 = w23818 ^ w23819;
	assign w9496 = w50110 ^ w50114;
	assign w9247 = w50115 ^ w50114;
	assign w45514 = ~w23928;
	assign w9501 = w45331 ^ w45514;
	assign w15867 = w46756 & w15881;
	assign w44030 = w15861 ^ w15867;
	assign w15773 = w15805 ^ w44030;
	assign w15816 = w46751 ^ w15773;
	assign w15851 = w15856 ^ w15816;
	assign w15850 = w15851 & w15852;
	assign w15849 = w15850 ^ w15858;
	assign w15835 = w15849 & w46756;
	assign w15768 = w15850 ^ w15867;
	assign w15848 = w15856 ^ w15850;
	assign w15847 = w15858 & w15848;
	assign w15845 = w15847 ^ w15855;
	assign w15763 = w15768 ^ w15864;
	assign w15826 = w15849 & w15881;
	assign w15769 = w15850 ^ w15814;
	assign w15811 = w44030 ^ w15796;
	assign w15857 = w15819 ^ w15811;
	assign w44035 = w15847 ^ w15865;
	assign w15839 = w44035 ^ w15817;
	assign w15828 = w15839 & w15880;
	assign w15837 = w15839 & w15876;
	assign w44034 = w15835 ^ w15837;
	assign w15806 = w46755 ^ w44035;
	assign w15846 = w15806 ^ w15769;
	assign w15827 = w15846 & w15877;
	assign w15854 = w15857 & w15855;
	assign w15853 = w15854 ^ w15816;
	assign w15823 = w15853 & w15879;
	assign w15765 = w15854 ^ w15866;
	assign w15761 = w15765 ^ w15801;
	assign w15844 = w15853 & w15845;
	assign w15832 = w15853 & w15872;
	assign w15767 = w15844 ^ w15868;
	assign w15759 = w15806 ^ w15767;
	assign w15766 = w15796 ^ w15759;
	assign w15842 = w15763 ^ w15766;
	assign w15829 = w15842 & w15874;
	assign w15820 = w15842 & w15883;
	assign w15764 = w46749 ^ w15761;
	assign w15841 = w15763 ^ w15764;
	assign w15831 = w15841 & w15873;
	assign w15822 = w15841 & w15884;
	assign w15786 = w15831 ^ w15820;
	assign w15762 = w15854 ^ w15810;
	assign w15782 = ~w15786;
	assign w15809 = w15844 ^ w15819;
	assign w15843 = w15809 ^ w15811;
	assign w15824 = w15843 & w15878;
	assign w15840 = w15809 ^ w15762;
	assign w15825 = w15840 & w15885;
	assign w15834 = w15840 & w15870;
	assign w15792 = w15834 ^ w15825;
	assign w15833 = w15843 & w15882;
	assign w15794 = w15832 ^ w15824;
	assign w15807 = w15825 ^ w15829;
	assign w15785 = ~w15807;
	assign w15784 = w15785 ^ w15823;
	assign w15780 = w15784 ^ w44034;
	assign w44033 = w15833 ^ w15834;
	assign w15783 = w15822 ^ w15780;
	assign w15887 = w15782 ^ w15783;
	assign w45326 = ~w15887;
	assign w9412 = w45326 ^ w33173;
	assign w15776 = w15832 ^ w15833;
	assign w15836 = w15846 & w15875;
	assign w15760 = w46751 ^ w15761;
	assign w15838 = w15759 ^ w15760;
	assign w15830 = w15838 & w15871;
	assign w15821 = w15838 & w15886;
	assign w15815 = w15830 ^ w44033;
	assign w15775 = w15831 ^ w15815;
	assign w15781 = w15826 ^ w15815;
	assign w15787 = w15830 ^ w15831;
	assign w44032 = w15821 ^ w15822;
	assign w15803 = w15827 ^ w44032;
	assign w15779 = w15803 ^ w15780;
	assign w15790 = w15794 ^ w44032;
	assign w15789 = w15785 ^ w15790;
	assign w15793 = w44034 ^ w15790;
	assign w15890 = w15792 ^ w15793;
	assign w15778 = ~w15781;
	assign w50056 = w15778 ^ w15779;
	assign w9281 = ~w50056;
	assign w9459 = w45340 ^ w9281;
	assign w9524 = w50049 ^ w50056;
	assign w9407 = ~w9524;
	assign w9418 = w9549 ^ w9407;
	assign w9405 = w9407 ^ w50045;
	assign w45328 = ~w15890;
	assign w9278 = w45340 ^ w45328;
	assign w9525 = w45766 ^ w45328;
	assign w15804 = w15828 ^ w15803;
	assign w15808 = w15836 ^ w15804;
	assign w15777 = w15835 ^ w15808;
	assign w15813 = w15837 ^ w15808;
	assign w50058 = w44033 ^ w15813;
	assign w9414 = w50058 ^ w50051;
	assign w15888 = w15813 ^ w15787;
	assign w45327 = ~w15888;
	assign w9410 = w45327 ^ w33174;
	assign w50057 = w15776 ^ w15777;
	assign w9280 = w50057 ^ w9281;
	assign w9272 = w50057 ^ w50050;
	assign w50059 = w15804 ^ w15775;
	assign w9486 = w50054 ^ w50059;
	assign w9420 = ~w9486;
	assign w9424 = w9420 ^ w45773;
	assign w15791 = w15830 ^ w15833;
	assign w15788 = ~w15791;
	assign w15889 = w15788 ^ w15789;
	assign w9274 = w15889 ^ w45341;
	assign w50055 = ~w15889;
	assign w9526 = w45773 ^ w50055;
	assign w26808 = w26830 & w26871;
	assign w26774 = w26819 ^ w26808;
	assign w26770 = ~w26774;
	assign w26875 = w26770 ^ w26771;
	assign w45600 = ~w26875;
	assign w23829 = w23825 ^ w23830;
	assign w23929 = w23828 ^ w23829;
	assign w45515 = ~w23929;
	assign w9508 = w45332 ^ w45515;
	assign w26803 = w26818 ^ w44494;
	assign w26769 = w26814 ^ w26803;
	assign w26763 = w26819 ^ w26803;
	assign w50085 = w26792 ^ w26763;
	assign w26766 = ~w26769;
	assign w50082 = w26766 ^ w26767;
	assign w45939 = ~w9134;
	assign w9122 = w45939 ^ w45369;
	assign w9117 = w45939 ^ w49910;
	assign w9120 = w9121 ^ w9122;
	assign w49821 = ~w9120;
	assign w49823 = w9116 ^ w9117;
	assign w46763 = w49821 ^ w968;
	assign w11597 = w46757 ^ w46763;
	assign w46761 = w49823 ^ w970;
	assign w11484 = w46761 ^ w46762;
	assign w11507 = w46763 ^ w46761;
	assign w11509 = w46762 ^ w11507;
	assign w11585 = w46758 ^ w11509;
	assign w11584 = w11514 ^ w11509;
	assign w11576 = w11591 & w11584;
	assign w11582 = w46759 ^ w11509;
	assign w11578 = w11597 & w11582;
	assign w11590 = w46763 ^ w11594;
	assign w11577 = w11594 & w11590;
	assign w8937 = w45939 ^ w49901;
	assign w9206 = w8937 ^ w8938;
	assign w49824 = w9206 ^ w9150;
	assign w46760 = w49824 ^ w971;
	assign w11510 = w46760 ^ w46758;
	assign w11470 = w11510 ^ w11508;
	assign w11586 = w11507 ^ w11470;
	assign w11573 = w11595 & w11586;
	assign w11469 = w11510 ^ w46759;
	assign w11593 = w46764 ^ w11469;
	assign w11579 = w46764 & w11593;
	assign w11512 = w11578 ^ w11508;
	assign w11524 = w46763 ^ w46762;
	assign w11589 = w11524 ^ w11591;
	assign w43854 = w11573 ^ w11576;
	assign w11486 = w11512 ^ w43854;
	assign w43853 = w11573 ^ w11579;
	assign w11523 = w43853 ^ w11508;
	assign w11598 = w46762 ^ w46760;
	assign w11583 = w11508 ^ w11598;
	assign w11574 = w11598 & w11583;
	assign w11526 = w11574 ^ w43854;
	assign w11482 = w11577 ^ w11526;
	assign w11564 = w46763 ^ w11482;
	assign w11596 = w46760 ^ w46757;
	assign w11575 = w11596 & w11585;
	assign w11483 = w11574 ^ w11575;
	assign w11530 = w11483 ^ w11484;
	assign w11529 = w11530 ^ w11512;
	assign w11588 = w11507 ^ w11596;
	assign w11511 = w11575 ^ w11509;
	assign w11570 = w11486 ^ w11511;
	assign w11571 = w11577 ^ w11529;
	assign w11587 = w46764 ^ w11588;
	assign w11580 = w11589 & w11587;
	assign w11531 = w11574 ^ w11580;
	assign w11569 = w11531 ^ w11523;
	assign w11592 = w11596 ^ w11524;
	assign w11581 = w11588 & w11592;
	assign w11513 = w11581 ^ w11510;
	assign w11517 = w11513 ^ w11511;
	assign w11485 = w11517 ^ w43853;
	assign w11528 = w46759 ^ w11485;
	assign w11522 = w46757 ^ w11517;
	assign w11572 = w11531 ^ w11522;
	assign w11568 = w11572 & w11571;
	assign w11563 = w11568 ^ w11528;
	assign w11562 = w11563 & w11564;
	assign w11561 = w11562 ^ w11570;
	assign w11538 = w11561 & w11593;
	assign w11481 = w11562 ^ w11526;
	assign w11480 = w11562 ^ w11579;
	assign w11475 = w11480 ^ w11576;
	assign w11547 = w11561 & w46764;
	assign w11567 = w11568 ^ w11570;
	assign w11566 = w11569 & w11567;
	assign w11474 = w11566 ^ w11522;
	assign w11477 = w11566 ^ w11578;
	assign w11473 = w11477 ^ w11513;
	assign w11476 = w46757 ^ w11473;
	assign w11553 = w11475 ^ w11476;
	assign w11534 = w11553 & w11596;
	assign w11472 = w46759 ^ w11473;
	assign w11565 = w11566 ^ w11528;
	assign w11535 = w11565 & w11591;
	assign w11544 = w11565 & w11584;
	assign w11560 = w11568 ^ w11562;
	assign w11559 = w11570 & w11560;
	assign w11557 = w11559 ^ w11567;
	assign w11556 = w11565 & w11557;
	assign w11479 = w11556 ^ w11580;
	assign w11521 = w11556 ^ w11531;
	assign w11552 = w11521 ^ w11474;
	assign w11555 = w11521 ^ w11523;
	assign w11536 = w11555 & w11590;
	assign w11506 = w11544 ^ w11536;
	assign w11546 = w11552 & w11582;
	assign w11545 = w11555 & w11594;
	assign w11488 = w11544 ^ w11545;
	assign w43855 = w11545 ^ w11546;
	assign w43857 = w11559 ^ w11577;
	assign w11518 = w46763 ^ w43857;
	assign w11558 = w11518 ^ w11481;
	assign w11548 = w11558 & w11587;
	assign w11539 = w11558 & w11589;
	assign w11471 = w11518 ^ w11479;
	assign w11478 = w11508 ^ w11471;
	assign w11554 = w11475 ^ w11478;
	assign w11541 = w11554 & w11586;
	assign w11532 = w11554 & w11595;
	assign w11550 = w11471 ^ w11472;
	assign w11533 = w11550 & w11598;
	assign w43528 = w11533 ^ w11534;
	assign w11502 = w11506 ^ w43528;
	assign w11515 = w11539 ^ w43528;
	assign w11542 = w11550 & w11583;
	assign w11527 = w11542 ^ w43855;
	assign w11493 = w11538 ^ w11527;
	assign w11503 = w11542 ^ w11545;
	assign w11500 = ~w11503;
	assign w11490 = ~w11493;
	assign w11543 = w11553 & w11585;
	assign w11498 = w11543 ^ w11532;
	assign w11487 = w11543 ^ w11527;
	assign w11499 = w11542 ^ w11543;
	assign w11494 = ~w11498;
	assign w11537 = w11552 & w11597;
	assign w11504 = w11546 ^ w11537;
	assign w11519 = w11537 ^ w11541;
	assign w11497 = ~w11519;
	assign w11501 = w11497 ^ w11502;
	assign w11601 = w11500 ^ w11501;
	assign w11496 = w11497 ^ w11535;
	assign w9237 = w11601 ^ w45337;
	assign w9570 = w9236 ^ w9237;
	assign w50069 = ~w11601;
	assign w9521 = w45336 ^ w50069;
	assign w11551 = w43857 ^ w11529;
	assign w11540 = w11551 & w11592;
	assign w11549 = w11551 & w11588;
	assign w43856 = w11547 ^ w11549;
	assign w11505 = w43856 ^ w11502;
	assign w11602 = w11504 ^ w11505;
	assign w11492 = w11496 ^ w43856;
	assign w11495 = w11534 ^ w11492;
	assign w11599 = w11494 ^ w11495;
	assign w11491 = w11515 ^ w11492;
	assign w50070 = w11490 ^ w11491;
	assign w9396 = w50070 ^ w45336;
	assign w9517 = w50065 ^ w50070;
	assign w9370 = ~w9517;
	assign w9368 = w9370 ^ w50078;
	assign w45231 = ~w11599;
	assign w9506 = w45334 ^ w45231;
	assign w9394 = w45231 ^ w50067;
	assign w9374 = w9506 ^ w9500;
	assign w45233 = ~w11602;
	assign w9522 = w45337 ^ w45233;
	assign w9367 = w9506 ^ w45686;
	assign w9365 = ~w9367;
	assign w11516 = w11540 ^ w11515;
	assign w50073 = w11516 ^ w11487;
	assign w9482 = w50068 ^ w50073;
	assign w11520 = w11548 ^ w11516;
	assign w11525 = w11549 ^ w11520;
	assign w11489 = w11547 ^ w11520;
	assign w50071 = w11488 ^ w11489;
	assign w11600 = w11525 ^ w11499;
	assign w9241 = ~w50071;
	assign w9240 = w9241 ^ w50065;
	assign w9569 = w9239 ^ w9240;
	assign w9514 = w50066 ^ w50071;
	assign w9378 = ~w9514;
	assign w9345 = w9482 ^ w45687;
	assign w45232 = ~w11600;
	assign w9364 = w45232 ^ w45231;
	assign w50072 = w43855 ^ w11525;
	assign w9510 = w50067 ^ w50072;
	assign w9243 = w50072 ^ w50066;
	assign w9568 = w9242 ^ w9243;
	assign w9352 = ~w9510;
	assign w45940 = ~w9140;
	assign w9064 = w45940 ^ w49863;
	assign w49739 = w9064 ^ w9065;
	assign w9085 = w45940 ^ w49846;
	assign w49728 = w9084 ^ w9085;
	assign w46845 = w49739 ^ w1077;
	assign w16332 = w46847 ^ w46845;
	assign w16294 = w16334 ^ w16332;
	assign w16410 = w16331 ^ w16294;
	assign w16407 = w16332 ^ w16422;
	assign w16398 = w16422 & w16407;
	assign w16421 = w46845 ^ w46851;
	assign w16402 = w16421 & w16406;
	assign w46856 = w49728 ^ w1066;
	assign w11778 = w46856 ^ w46854;
	assign w11864 = w46856 ^ w46853;
	assign w11866 = w46858 ^ w46856;
	assign w11851 = w11776 ^ w11866;
	assign w11842 = w11866 & w11851;
	assign w11738 = w11778 ^ w11776;
	assign w11737 = w11778 ^ w46855;
	assign w11861 = w46860 ^ w11737;
	assign w11847 = w46860 & w11861;
	assign w8928 = w45940 ^ w45241;
	assign w9210 = w8928 ^ w8929;
	assign w49725 = w9210 ^ w9202;
	assign w46859 = w49725 ^ w1063;
	assign w11858 = w46859 ^ w11862;
	assign w11775 = w46859 ^ w46857;
	assign w11777 = w46858 ^ w11775;
	assign w11852 = w11782 ^ w11777;
	assign w11853 = w46854 ^ w11777;
	assign w11850 = w46855 ^ w11777;
	assign w11856 = w11775 ^ w11864;
	assign w11855 = w46860 ^ w11856;
	assign w11792 = w46859 ^ w46858;
	assign w11857 = w11792 ^ w11859;
	assign w11860 = w11864 ^ w11792;
	assign w11844 = w11859 & w11852;
	assign w11865 = w46853 ^ w46859;
	assign w11848 = w11857 & w11855;
	assign w11799 = w11842 ^ w11848;
	assign w11849 = w11856 & w11860;
	assign w11781 = w11849 ^ w11778;
	assign w11854 = w11775 ^ w11738;
	assign w11846 = w11865 & w11850;
	assign w11780 = w11846 ^ w11776;
	assign w11845 = w11862 & w11858;
	assign w11843 = w11864 & w11853;
	assign w11779 = w11843 ^ w11777;
	assign w11785 = w11781 ^ w11779;
	assign w11751 = w11842 ^ w11843;
	assign w11790 = w46853 ^ w11785;
	assign w11840 = w11799 ^ w11790;
	assign w11798 = w11751 ^ w11752;
	assign w11797 = w11798 ^ w11780;
	assign w11839 = w11845 ^ w11797;
	assign w11836 = w11840 & w11839;
	assign w16419 = w46845 ^ w46850;
	assign w16397 = w16419 & w16410;
	assign w44053 = w16397 ^ w16403;
	assign w16336 = w16402 ^ w16332;
	assign w16420 = w46848 ^ w46845;
	assign w16399 = w16420 & w16409;
	assign w16307 = w16398 ^ w16399;
	assign w16416 = w16420 ^ w16348;
	assign w16354 = w16307 ^ w16308;
	assign w16412 = w16331 ^ w16420;
	assign w16405 = w16412 & w16416;
	assign w16353 = w16354 ^ w16336;
	assign w16395 = w16401 ^ w16353;
	assign w16411 = w46852 ^ w16412;
	assign w16335 = w16399 ^ w16333;
	assign w16337 = w16405 ^ w16334;
	assign w11841 = w11863 & w11854;
	assign w43864 = w11841 ^ w11847;
	assign w11791 = w43864 ^ w11776;
	assign w11837 = w11799 ^ w11791;
	assign w11753 = w11785 ^ w43864;
	assign w11796 = w46855 ^ w11753;
	assign w11831 = w11836 ^ w11796;
	assign w43865 = w11841 ^ w11844;
	assign w11794 = w11842 ^ w43865;
	assign w11750 = w11845 ^ w11794;
	assign w11832 = w46859 ^ w11750;
	assign w11830 = w11831 & w11832;
	assign w11828 = w11836 ^ w11830;
	assign w11748 = w11830 ^ w11847;
	assign w11743 = w11748 ^ w11844;
	assign w11749 = w11830 ^ w11794;
	assign w11754 = w11780 ^ w43865;
	assign w11838 = w11754 ^ w11779;
	assign w11829 = w11830 ^ w11838;
	assign w11835 = w11836 ^ w11838;
	assign w11834 = w11837 & w11835;
	assign w11742 = w11834 ^ w11790;
	assign w11833 = w11834 ^ w11796;
	assign w11745 = w11834 ^ w11846;
	assign w11827 = w11838 & w11828;
	assign w11825 = w11827 ^ w11835;
	assign w11824 = w11833 & w11825;
	assign w11789 = w11824 ^ w11799;
	assign w11823 = w11789 ^ w11791;
	assign w11747 = w11824 ^ w11848;
	assign w11741 = w11745 ^ w11781;
	assign w11740 = w46855 ^ w11741;
	assign w11815 = w11829 & w46860;
	assign w11744 = w46853 ^ w11741;
	assign w11821 = w11743 ^ w11744;
	assign w11811 = w11821 & w11853;
	assign w11813 = w11823 & w11862;
	assign w11812 = w11833 & w11852;
	assign w11756 = w11812 ^ w11813;
	assign w11820 = w11789 ^ w11742;
	assign w11814 = w11820 & w11850;
	assign w11803 = w11833 & w11859;
	assign w11804 = w11823 & w11858;
	assign w11774 = w11812 ^ w11804;
	assign w11806 = w11829 & w11861;
	assign w11805 = w11820 & w11865;
	assign w11772 = w11814 ^ w11805;
	assign w11802 = w11821 & w11864;
	assign w43866 = w11813 ^ w11814;
	assign w43868 = w11827 ^ w11845;
	assign w11786 = w46859 ^ w43868;
	assign w11826 = w11786 ^ w11749;
	assign w11807 = w11826 & w11857;
	assign w11816 = w11826 & w11855;
	assign w11739 = w11786 ^ w11747;
	assign w11818 = w11739 ^ w11740;
	assign w11801 = w11818 & w11866;
	assign w43529 = w11801 ^ w11802;
	assign w11770 = w11774 ^ w43529;
	assign w11746 = w11776 ^ w11739;
	assign w11822 = w11743 ^ w11746;
	assign w11800 = w11822 & w11863;
	assign w11766 = w11811 ^ w11800;
	assign w11762 = ~w11766;
	assign w11809 = w11822 & w11854;
	assign w11787 = w11805 ^ w11809;
	assign w11765 = ~w11787;
	assign w11764 = w11765 ^ w11803;
	assign w11769 = w11765 ^ w11770;
	assign w11810 = w11818 & w11851;
	assign w11771 = w11810 ^ w11813;
	assign w11767 = w11810 ^ w11811;
	assign w11768 = ~w11771;
	assign w11869 = w11768 ^ w11769;
	assign w50086 = ~w11869;
	assign w9545 = w45594 ^ w50086;
	assign w9313 = w45598 ^ w11869;
	assign w9256 = w11869 ^ w45595;
	assign w11819 = w43868 ^ w11797;
	assign w11808 = w11819 & w11860;
	assign w11783 = w11807 ^ w43529;
	assign w11784 = w11808 ^ w11783;
	assign w11788 = w11816 ^ w11784;
	assign w11757 = w11815 ^ w11788;
	assign w50088 = w11756 ^ w11757;
	assign w9531 = w50083 ^ w50088;
	assign w9260 = ~w50088;
	assign w9270 = w50094 ^ w9260;
	assign w9259 = w9260 ^ w50082;
	assign w9298 = ~w9531;
	assign w11795 = w11810 ^ w43866;
	assign w11755 = w11811 ^ w11795;
	assign w50092 = w11784 ^ w11755;
	assign w9331 = w50092 ^ w45601;
	assign w11761 = w11806 ^ w11795;
	assign w11758 = ~w11761;
	assign w9487 = w50092 ^ w50096;
	assign w9483 = w50085 ^ w50092;
	assign w9268 = ~w9487;
	assign w11817 = w11819 & w11856;
	assign w43867 = w11815 ^ w11817;
	assign w11773 = w43867 ^ w11770;
	assign w11870 = w11772 ^ w11773;
	assign w11760 = w11764 ^ w43867;
	assign w11759 = w11783 ^ w11760;
	assign w11763 = w11802 ^ w11760;
	assign w11867 = w11762 ^ w11763;
	assign w9308 = w45604 ^ w11867;
	assign w9339 = w11867 ^ w50084;
	assign w50087 = w11758 ^ w11759;
	assign w9267 = ~w50087;
	assign w9266 = w50093 ^ w9267;
	assign w9538 = w50082 ^ w50087;
	assign w9314 = ~w9538;
	assign w50090 = ~w11867;
	assign w9516 = w45600 ^ w50090;
	assign w11793 = w11817 ^ w11788;
	assign w11868 = w11793 ^ w11767;
	assign w9334 = w11868 ^ w45600;
	assign w9306 = w45605 ^ w11868;
	assign w50089 = w43866 ^ w11793;
	assign w9311 = w50095 ^ w50089;
	assign w50091 = ~w11868;
	assign w9509 = w45601 ^ w50091;
	assign w9523 = w50084 ^ w50089;
	assign w9295 = ~w9523;
	assign w9262 = w50089 ^ w50083;
	assign w45234 = ~w11870;
	assign w9264 = w45599 ^ w45234;
	assign w9546 = w45595 ^ w45234;
	assign w16347 = w44053 ^ w16332;
	assign w16341 = w16337 ^ w16335;
	assign w16309 = w16341 ^ w44053;
	assign w16352 = w46847 ^ w16309;
	assign w16346 = w46845 ^ w16341;
	assign w16415 = w16332 ^ w16338;
	assign w16400 = w16415 & w16408;
	assign w16413 = w16348 ^ w16415;
	assign w16404 = w16413 & w16411;
	assign w44054 = w16397 ^ w16400;
	assign w16310 = w16336 ^ w44054;
	assign w16394 = w16310 ^ w16335;
	assign w16350 = w16398 ^ w44054;
	assign w16306 = w16401 ^ w16350;
	assign w16388 = w46851 ^ w16306;
	assign w9342 = w9267 ^ w45594;
	assign w9315 = w9546 ^ w9487;
	assign w16355 = w16398 ^ w16404;
	assign w16396 = w16355 ^ w16346;
	assign w16392 = w16396 & w16395;
	assign w16387 = w16392 ^ w16352;
	assign w16386 = w16387 & w16388;
	assign w16304 = w16386 ^ w16403;
	assign w16299 = w16304 ^ w16400;
	assign w16305 = w16386 ^ w16350;
	assign w16385 = w16386 ^ w16394;
	assign w16371 = w16385 & w46852;
	assign w16362 = w16385 & w16417;
	assign w16384 = w16392 ^ w16386;
	assign w16383 = w16394 & w16384;
	assign w44057 = w16383 ^ w16401;
	assign w16342 = w46851 ^ w44057;
	assign w16382 = w16342 ^ w16305;
	assign w16363 = w16382 & w16413;
	assign w16372 = w16382 & w16411;
	assign w16375 = w44057 ^ w16353;
	assign w16364 = w16375 & w16416;
	assign w16373 = w16375 & w16412;
	assign w44056 = w16371 ^ w16373;
	assign w16391 = w16392 ^ w16394;
	assign w16381 = w16383 ^ w16391;
	assign w16393 = w16355 ^ w16347;
	assign w16390 = w16393 & w16391;
	assign w16298 = w16390 ^ w16346;
	assign w16301 = w16390 ^ w16402;
	assign w16297 = w16301 ^ w16337;
	assign w16296 = w46847 ^ w16297;
	assign w16300 = w46845 ^ w16297;
	assign w16377 = w16299 ^ w16300;
	assign w16358 = w16377 & w16420;
	assign w16367 = w16377 & w16409;
	assign w45896 = ~w9483;
	assign w9322 = w45896 ^ w50084;
	assign w9324 = w45896 ^ w50083;
	assign w9328 = w45896 ^ w45594;
	assign w16389 = w16390 ^ w16352;
	assign w16368 = w16389 & w16408;
	assign w16380 = w16389 & w16381;
	assign w16345 = w16380 ^ w16355;
	assign w16303 = w16380 ^ w16404;
	assign w16295 = w16342 ^ w16303;
	assign w16376 = w16345 ^ w16298;
	assign w16374 = w16295 ^ w16296;
	assign w16302 = w16332 ^ w16295;
	assign w16378 = w16299 ^ w16302;
	assign w16379 = w16345 ^ w16347;
	assign w16365 = w16378 & w16410;
	assign w16366 = w16374 & w16407;
	assign w16323 = w16366 ^ w16367;
	assign w16370 = w16376 & w16406;
	assign w16361 = w16376 & w16421;
	assign w16343 = w16361 ^ w16365;
	assign w16321 = ~w16343;
	assign w16356 = w16378 & w16419;
	assign w16322 = w16367 ^ w16356;
	assign w16318 = ~w16322;
	assign w16369 = w16379 & w16418;
	assign w16312 = w16368 ^ w16369;
	assign w16357 = w16374 & w16422;
	assign w16360 = w16379 & w16414;
	assign w16330 = w16368 ^ w16360;
	assign w16359 = w16389 & w16415;
	assign w16320 = w16321 ^ w16359;
	assign w16316 = w16320 ^ w44056;
	assign w16319 = w16358 ^ w16316;
	assign w16423 = w16318 ^ w16319;
	assign w43544 = w16357 ^ w16358;
	assign w16339 = w16363 ^ w43544;
	assign w16315 = w16339 ^ w16316;
	assign w16340 = w16364 ^ w16339;
	assign w16344 = w16372 ^ w16340;
	assign w16313 = w16371 ^ w16344;
	assign w50075 = w16312 ^ w16313;
	assign w9253 = w50075 ^ w9241;
	assign w9507 = w50075 ^ w50079;
	assign w9349 = w9352 ^ w9507;
	assign w16349 = w16373 ^ w16344;
	assign w16424 = w16349 ^ w16323;
	assign w9379 = w9370 ^ w9507;
	assign w49952 = w9569 ^ w9507;
	assign w46705 = w49952 ^ w1153;
	assign w44055 = w16369 ^ w16370;
	assign w50076 = w44055 ^ w16349;
	assign w9351 = ~w50076;
	assign w9366 = w9351 ^ w50072;
	assign w9502 = w50076 ^ w50080;
	assign w9348 = w9506 ^ w9502;
	assign w49953 = w9568 ^ w9502;
	assign w46704 = w49953 ^ w1154;
	assign w9376 = w9378 ^ w9502;
	assign w49970 = w9365 ^ w9366;
	assign w46687 = w49970 ^ w1171;
	assign w45342 = ~w16423;
	assign w9363 = w9500 ^ w45342;
	assign w49978 = w45342 ^ w9348;
	assign w46679 = w49978 ^ w1179;
	assign w9497 = w45342 ^ w45686;
	assign w9393 = w9497 ^ w50080;
	assign w49954 = w9393 ^ w9394;
	assign w46703 = w49954 ^ w1155;
	assign w9375 = w9510 ^ w9497;
	assign w49962 = w45334 ^ w9375;
	assign w46695 = w49962 ^ w1163;
	assign w49971 = w9363 ^ w9364;
	assign w46686 = w49971 ^ w1172;
	assign w45343 = ~w16424;
	assign w49963 = w45343 ^ w9374;
	assign w46694 = w49963 ^ w1164;
	assign w9499 = w45232 ^ w45343;
	assign w9362 = w9499 ^ w9482;
	assign w9347 = w9499 ^ w9497;
	assign w9391 = w9499 ^ w45687;
	assign w49979 = w45335 ^ w9347;
	assign w46678 = w49979 ^ w1180;
	assign w49972 = w50081 ^ w9362;
	assign w46685 = w49972 ^ w1173;
	assign w15394 = w46687 ^ w46685;
	assign w16351 = w16366 ^ w44055;
	assign w16311 = w16367 ^ w16351;
	assign w50077 = w16340 ^ w16311;
	assign w16317 = w16362 ^ w16351;
	assign w16314 = ~w16317;
	assign w50074 = w16314 ^ w16315;
	assign w9251 = w50074 ^ w50070;
	assign w9346 = w50077 ^ w45343;
	assign w49980 = w9345 ^ w9346;
	assign w46677 = w49980 ^ w1181;
	assign w29598 = w46679 ^ w46677;
	assign w9489 = w50073 ^ w50077;
	assign w9254 = ~w9489;
	assign w9252 = w9254 ^ w50080;
	assign w9248 = w9489 ^ w45688;
	assign w9481 = w50077 ^ w50081;
	assign w9361 = w9522 ^ w9481;
	assign w9357 = w9481 ^ w50075;
	assign w9372 = w9481 ^ w45232;
	assign w49964 = w9372 ^ w9373;
	assign w46693 = w49964 ^ w1165;
	assign w32948 = w46695 ^ w46693;
	assign w9390 = w9500 ^ w9481;
	assign w49956 = w50073 ^ w9390;
	assign w46701 = w49956 ^ w1157;
	assign w15616 = w46704 ^ w46701;
	assign w15528 = w46703 ^ w46701;
	assign w9250 = w9489 ^ w50079;
	assign w9564 = w9250 ^ w9251;
	assign w49968 = w9564 ^ w9514;
	assign w46689 = w49968 ^ w1169;
	assign w9512 = w50074 ^ w50078;
	assign w9381 = w9521 ^ w9512;
	assign w9395 = w9512 ^ w45688;
	assign w49951 = w9395 ^ w9396;
	assign w46706 = w49951 ^ w1152;
	assign w15615 = w46701 ^ w46706;
	assign w15504 = w46705 ^ w46706;
	assign w15618 = w46706 ^ w46704;
	assign w49959 = w50065 ^ w9381;
	assign w46698 = w49959 ^ w1160;
	assign w33035 = w46693 ^ w46698;
	assign w9371 = w9522 ^ w9489;
	assign w49965 = w45689 ^ w9371;
	assign w46692 = w49965 ^ w1166;
	assign w15400 = w46692 ^ w46686;
	assign w15480 = w46687 ^ w15400;
	assign w15477 = w15394 ^ w15400;
	assign w9356 = w9514 ^ w9512;
	assign w49976 = w9356 ^ w9357;
	assign w46681 = w49976 ^ w1177;
	assign w9350 = w9481 ^ w9351;
	assign w49977 = w9349 ^ w9350;
	assign w46680 = w49977 ^ w1178;
	assign w29686 = w46680 ^ w46677;
	assign w29600 = w46680 ^ w46678;
	assign w29559 = w29600 ^ w46679;
	assign w29560 = w29600 ^ w29598;
	assign w9563 = w9252 ^ w9253;
	assign w49969 = w9563 ^ w9510;
	assign w46688 = w49969 ^ w1170;
	assign w15396 = w46688 ^ w46686;
	assign w15355 = w15396 ^ w46687;
	assign w15479 = w46692 ^ w15355;
	assign w15465 = w46692 & w15479;
	assign w15356 = w15396 ^ w15394;
	assign w15482 = w46688 ^ w46685;
	assign w16328 = w16370 ^ w16361;
	assign w16326 = w16330 ^ w43544;
	assign w16329 = w44056 ^ w16326;
	assign w16426 = w16328 ^ w16329;
	assign w45345 = ~w16426;
	assign w49973 = w45345 ^ w9361;
	assign w46684 = w49973 ^ w1174;
	assign w29683 = w46684 ^ w29559;
	assign w29604 = w46684 ^ w46678;
	assign w9249 = w45345 ^ w45233;
	assign w9565 = w9248 ^ w9249;
	assign w29684 = w46679 ^ w29604;
	assign w29681 = w29598 ^ w29604;
	assign w9519 = w45345 ^ w45689;
	assign w9359 = w9521 ^ w9519;
	assign w9397 = w9519 ^ w9491;
	assign w49949 = w45233 ^ w9397;
	assign w46708 = w49949 ^ w1150;
	assign w29669 = w46684 & w29683;
	assign w9385 = w9519 ^ w9482;
	assign w49957 = w45337 ^ w9385;
	assign w46700 = w49957 ^ w1158;
	assign w32954 = w46700 ^ w46694;
	assign w33031 = w32948 ^ w32954;
	assign w33034 = w46695 ^ w32954;
	assign w49966 = w9565 ^ w9521;
	assign w46691 = w49966 ^ w1167;
	assign w15393 = w46691 ^ w46689;
	assign w15472 = w15393 ^ w15356;
	assign w15474 = w15393 ^ w15482;
	assign w15473 = w46692 ^ w15474;
	assign w15476 = w46691 ^ w15480;
	assign w15463 = w15480 & w15476;
	assign w15483 = w46685 ^ w46691;
	assign w16325 = w16321 ^ w16326;
	assign w15603 = w15528 ^ w15618;
	assign w15594 = w15618 & w15603;
	assign w49955 = w9391 ^ w9392;
	assign w46702 = w49955 ^ w1156;
	assign w15534 = w46708 ^ w46702;
	assign w15611 = w15528 ^ w15534;
	assign w15614 = w46703 ^ w15534;
	assign w15530 = w46704 ^ w46702;
	assign w15489 = w15530 ^ w46703;
	assign w15613 = w46708 ^ w15489;
	assign w15599 = w46708 & w15613;
	assign w15490 = w15530 ^ w15528;
	assign w16327 = w16366 ^ w16369;
	assign w16324 = ~w16327;
	assign w16425 = w16324 ^ w16325;
	assign w45344 = ~w16425;
	assign w9369 = w45344 ^ w11601;
	assign w9360 = w9481 ^ w45344;
	assign w9515 = w45344 ^ w45688;
	assign w9383 = w9522 ^ w9515;
	assign w49950 = w9570 ^ w9515;
	assign w46707 = w49950 ^ w1151;
	assign w15610 = w46707 ^ w15614;
	assign w15597 = w15614 & w15610;
	assign w15527 = w46707 ^ w46705;
	assign w15608 = w15527 ^ w15616;
	assign w15607 = w46708 ^ w15608;
	assign w15606 = w15527 ^ w15490;
	assign w15593 = w15615 & w15606;
	assign w15529 = w46706 ^ w15527;
	assign w15544 = w46707 ^ w46706;
	assign w15612 = w15616 ^ w15544;
	assign w15601 = w15608 & w15612;
	assign w15533 = w15601 ^ w15530;
	assign w15602 = w46703 ^ w15529;
	assign w15617 = w46701 ^ w46707;
	assign w15598 = w15617 & w15602;
	assign w15609 = w15544 ^ w15611;
	assign w15532 = w15598 ^ w15528;
	assign w44020 = w15593 ^ w15599;
	assign w15543 = w44020 ^ w15528;
	assign w49967 = w9368 ^ w9369;
	assign w46690 = w49967 ^ w1168;
	assign w15395 = w46690 ^ w15393;
	assign w15471 = w46686 ^ w15395;
	assign w15461 = w15482 & w15471;
	assign w15397 = w15461 ^ w15395;
	assign w15481 = w46685 ^ w46690;
	assign w15459 = w15481 & w15472;
	assign w15468 = w46687 ^ w15395;
	assign w15464 = w15483 & w15468;
	assign w15398 = w15464 ^ w15394;
	assign w44017 = w15459 ^ w15465;
	assign w15409 = w44017 ^ w15394;
	assign w15484 = w46690 ^ w46688;
	assign w15469 = w15394 ^ w15484;
	assign w15460 = w15484 & w15469;
	assign w15369 = w15460 ^ w15461;
	assign w15410 = w46691 ^ w46690;
	assign w15475 = w15410 ^ w15477;
	assign w15478 = w15482 ^ w15410;
	assign w15467 = w15474 & w15478;
	assign w15399 = w15467 ^ w15396;
	assign w15466 = w15475 & w15473;
	assign w15417 = w15460 ^ w15466;
	assign w15455 = w15417 ^ w15409;
	assign w15470 = w15400 ^ w15395;
	assign w15462 = w15477 & w15470;
	assign w44014 = w15459 ^ w15462;
	assign w15372 = w15398 ^ w44014;
	assign w15456 = w15372 ^ w15397;
	assign w15412 = w15460 ^ w44014;
	assign w15368 = w15463 ^ w15412;
	assign w15450 = w46691 ^ w15368;
	assign w49974 = w9359 ^ w9360;
	assign w46683 = w49974 ^ w1175;
	assign w29687 = w46677 ^ w46683;
	assign w29680 = w46683 ^ w29684;
	assign w29667 = w29684 & w29680;
	assign w9358 = w9517 ^ w9515;
	assign w49975 = w50074 ^ w9358;
	assign w46682 = w49975 ^ w1176;
	assign w29685 = w46677 ^ w46682;
	assign w29688 = w46682 ^ w46680;
	assign w29673 = w29598 ^ w29688;
	assign w29664 = w29688 & w29673;
	assign w29574 = w46681 ^ w46682;
	assign w15600 = w15609 & w15607;
	assign w15403 = w15399 ^ w15397;
	assign w15408 = w46685 ^ w15403;
	assign w15458 = w15417 ^ w15408;
	assign w15371 = w15403 ^ w44017;
	assign w15414 = w46687 ^ w15371;
	assign w15551 = w15594 ^ w15600;
	assign w15589 = w15551 ^ w15543;
	assign w15605 = w46702 ^ w15529;
	assign w15595 = w15616 & w15605;
	assign w15503 = w15594 ^ w15595;
	assign w15550 = w15503 ^ w15504;
	assign w15549 = w15550 ^ w15532;
	assign w15591 = w15597 ^ w15549;
	assign w15531 = w15595 ^ w15529;
	assign w15537 = w15533 ^ w15531;
	assign w15542 = w46701 ^ w15537;
	assign w15592 = w15551 ^ w15542;
	assign w15588 = w15592 & w15591;
	assign w29597 = w46683 ^ w46681;
	assign w29678 = w29597 ^ w29686;
	assign w29676 = w29597 ^ w29560;
	assign w29677 = w46684 ^ w29678;
	assign w29663 = w29685 & w29676;
	assign w44612 = w29663 ^ w29669;
	assign w29613 = w44612 ^ w29598;
	assign w29614 = w46683 ^ w46682;
	assign w29682 = w29686 ^ w29614;
	assign w29671 = w29678 & w29682;
	assign w29603 = w29671 ^ w29600;
	assign w15505 = w15537 ^ w44020;
	assign w15548 = w46703 ^ w15505;
	assign w15583 = w15588 ^ w15548;
	assign w15604 = w15534 ^ w15529;
	assign w15596 = w15611 & w15604;
	assign w44021 = w15593 ^ w15596;
	assign w15546 = w15594 ^ w44021;
	assign w15506 = w15532 ^ w44021;
	assign w15590 = w15506 ^ w15531;
	assign w15587 = w15588 ^ w15590;
	assign w15586 = w15589 & w15587;
	assign w15585 = w15586 ^ w15548;
	assign w15564 = w15585 & w15604;
	assign w15497 = w15586 ^ w15598;
	assign w15494 = w15586 ^ w15542;
	assign w15555 = w15585 & w15611;
	assign w15493 = w15497 ^ w15533;
	assign w15496 = w46701 ^ w15493;
	assign w15492 = w46703 ^ w15493;
	assign w29679 = w29614 ^ w29681;
	assign w29670 = w29679 & w29677;
	assign w29621 = w29664 ^ w29670;
	assign w29659 = w29621 ^ w29613;
	assign w15502 = w15597 ^ w15546;
	assign w15584 = w46707 ^ w15502;
	assign w15582 = w15583 & w15584;
	assign w15580 = w15588 ^ w15582;
	assign w15579 = w15590 & w15580;
	assign w15577 = w15579 ^ w15587;
	assign w15501 = w15582 ^ w15546;
	assign w15500 = w15582 ^ w15599;
	assign w15495 = w15500 ^ w15596;
	assign w15573 = w15495 ^ w15496;
	assign w15563 = w15573 & w15605;
	assign w15554 = w15573 & w15616;
	assign w44024 = w15579 ^ w15597;
	assign w15538 = w46707 ^ w44024;
	assign w15578 = w15538 ^ w15501;
	assign w15559 = w15578 & w15609;
	assign w15568 = w15578 & w15607;
	assign w15571 = w44024 ^ w15549;
	assign w15569 = w15571 & w15608;
	assign w15576 = w15585 & w15577;
	assign w15541 = w15576 ^ w15551;
	assign w15572 = w15541 ^ w15494;
	assign w15575 = w15541 ^ w15543;
	assign w15565 = w15575 & w15614;
	assign w15556 = w15575 & w15610;
	assign w15526 = w15564 ^ w15556;
	assign w15508 = w15564 ^ w15565;
	assign w15499 = w15576 ^ w15600;
	assign w15491 = w15538 ^ w15499;
	assign w15498 = w15528 ^ w15491;
	assign w15570 = w15491 ^ w15492;
	assign w15562 = w15570 & w15603;
	assign w15519 = w15562 ^ w15563;
	assign w15574 = w15495 ^ w15498;
	assign w15552 = w15574 & w15615;
	assign w15518 = w15563 ^ w15552;
	assign w15561 = w15574 & w15606;
	assign w15523 = w15562 ^ w15565;
	assign w15520 = ~w15523;
	assign w15514 = ~w15518;
	assign w15553 = w15570 & w15618;
	assign w43541 = w15553 ^ w15554;
	assign w15535 = w15559 ^ w43541;
	assign w15522 = w15526 ^ w43541;
	assign w15560 = w15571 & w15612;
	assign w15536 = w15560 ^ w15535;
	assign w15540 = w15568 ^ w15536;
	assign w15545 = w15569 ^ w15540;
	assign w15620 = w15545 ^ w15519;
	assign w45325 = ~w15620;
	assign w15566 = w15572 & w15602;
	assign w44022 = w15565 ^ w15566;
	assign w15547 = w15562 ^ w44022;
	assign w15507 = w15563 ^ w15547;
	assign w50249 = w15536 ^ w15507;
	assign w50248 = w44022 ^ w15545;
	assign w29599 = w46682 ^ w29597;
	assign w29674 = w29604 ^ w29599;
	assign w29666 = w29681 & w29674;
	assign w44609 = w29663 ^ w29666;
	assign w29616 = w29664 ^ w44609;
	assign w29675 = w46678 ^ w29599;
	assign w29665 = w29686 & w29675;
	assign w29573 = w29664 ^ w29665;
	assign w29601 = w29665 ^ w29599;
	assign w29607 = w29603 ^ w29601;
	assign w29575 = w29607 ^ w44612;
	assign w29612 = w46677 ^ w29607;
	assign w29618 = w46679 ^ w29575;
	assign w29662 = w29621 ^ w29612;
	assign w29672 = w46679 ^ w29599;
	assign w29668 = w29687 & w29672;
	assign w29602 = w29668 ^ w29598;
	assign w29576 = w29602 ^ w44609;
	assign w29660 = w29576 ^ w29601;
	assign w29620 = w29573 ^ w29574;
	assign w29619 = w29620 ^ w29602;
	assign w29661 = w29667 ^ w29619;
	assign w15581 = w15582 ^ w15590;
	assign w15567 = w15581 & w46708;
	assign w15558 = w15581 & w15613;
	assign w15513 = w15558 ^ w15547;
	assign w15509 = w15567 ^ w15540;
	assign w50247 = w15508 ^ w15509;
	assign w15510 = ~w15513;
	assign w44023 = w15567 ^ w15569;
	assign w15525 = w44023 ^ w15522;
	assign w29658 = w29662 & w29661;
	assign w29657 = w29658 ^ w29660;
	assign w29656 = w29659 & w29657;
	assign w29655 = w29656 ^ w29618;
	assign w29567 = w29656 ^ w29668;
	assign w29563 = w29567 ^ w29603;
	assign w29625 = w29655 & w29681;
	assign w29653 = w29658 ^ w29618;
	assign w29634 = w29655 & w29674;
	assign w29566 = w46677 ^ w29563;
	assign w29564 = w29656 ^ w29612;
	assign w15557 = w15572 & w15617;
	assign w15539 = w15557 ^ w15561;
	assign w15524 = w15566 ^ w15557;
	assign w15622 = w15524 ^ w15525;
	assign w45319 = ~w15622;
	assign w15517 = ~w15539;
	assign w15521 = w15517 ^ w15522;
	assign w15516 = w15517 ^ w15555;
	assign w15621 = w15520 ^ w15521;
	assign w15512 = w15516 ^ w44023;
	assign w15515 = w15554 ^ w15512;
	assign w15511 = w15535 ^ w15512;
	assign w15619 = w15514 ^ w15515;
	assign w50246 = w15510 ^ w15511;
	assign w45318 = ~w15621;
	assign w45324 = ~w15619;
	assign w15370 = w46689 ^ w46690;
	assign w15416 = w15369 ^ w15370;
	assign w15415 = w15416 ^ w15398;
	assign w15457 = w15463 ^ w15415;
	assign w15454 = w15458 & w15457;
	assign w15449 = w15454 ^ w15414;
	assign w15453 = w15454 ^ w15456;
	assign w15452 = w15455 & w15453;
	assign w15451 = w15452 ^ w15414;
	assign w15421 = w15451 & w15477;
	assign w15430 = w15451 & w15470;
	assign w15363 = w15452 ^ w15464;
	assign w15359 = w15363 ^ w15399;
	assign w15360 = w15452 ^ w15408;
	assign w15362 = w46685 ^ w15359;
	assign w15448 = w15449 & w15450;
	assign w15447 = w15448 ^ w15456;
	assign w15446 = w15454 ^ w15448;
	assign w15433 = w15447 & w46692;
	assign w15367 = w15448 ^ w15412;
	assign w15445 = w15456 & w15446;
	assign w44016 = w15445 ^ w15463;
	assign w15437 = w44016 ^ w15415;
	assign w15426 = w15437 & w15478;
	assign w15435 = w15437 & w15474;
	assign w15404 = w46691 ^ w44016;
	assign w15444 = w15404 ^ w15367;
	assign w15434 = w15444 & w15473;
	assign w15425 = w15444 & w15475;
	assign w44019 = w15433 ^ w15435;
	assign w15424 = w15447 & w15479;
	assign w15443 = w15445 ^ w15453;
	assign w15442 = w15451 & w15443;
	assign w15365 = w15442 ^ w15466;
	assign w15357 = w15404 ^ w15365;
	assign w15407 = w15442 ^ w15417;
	assign w15438 = w15407 ^ w15360;
	assign w15441 = w15407 ^ w15409;
	assign w15423 = w15438 & w15483;
	assign w15432 = w15438 & w15468;
	assign w15431 = w15441 & w15480;
	assign w15374 = w15430 ^ w15431;
	assign w15390 = w15432 ^ w15423;
	assign w15364 = w15394 ^ w15357;
	assign w44018 = w15431 ^ w15432;
	assign w15422 = w15441 & w15476;
	assign w15392 = w15430 ^ w15422;
	assign w15366 = w15448 ^ w15465;
	assign w15361 = w15366 ^ w15462;
	assign w15440 = w15361 ^ w15364;
	assign w15427 = w15440 & w15472;
	assign w15405 = w15423 ^ w15427;
	assign w15383 = ~w15405;
	assign w15382 = w15383 ^ w15421;
	assign w15378 = w15382 ^ w44019;
	assign w15439 = w15361 ^ w15362;
	assign w15429 = w15439 & w15471;
	assign w15420 = w15439 & w15482;
	assign w15381 = w15420 ^ w15378;
	assign w15418 = w15440 & w15481;
	assign w15384 = w15429 ^ w15418;
	assign w15380 = ~w15384;
	assign w15485 = w15380 ^ w15381;
	assign w45320 = ~w15485;
	assign w15358 = w46687 ^ w15359;
	assign w15436 = w15357 ^ w15358;
	assign w15428 = w15436 & w15469;
	assign w15385 = w15428 ^ w15429;
	assign w15389 = w15428 ^ w15431;
	assign w15386 = ~w15389;
	assign w15413 = w15428 ^ w44018;
	assign w15373 = w15429 ^ w15413;
	assign w15379 = w15424 ^ w15413;
	assign w15376 = ~w15379;
	assign w15419 = w15436 & w15484;
	assign w44015 = w15419 ^ w15420;
	assign w15401 = w15425 ^ w44015;
	assign w15402 = w15426 ^ w15401;
	assign w15406 = w15434 ^ w15402;
	assign w15375 = w15433 ^ w15406;
	assign w15411 = w15435 ^ w15406;
	assign w50296 = w44018 ^ w15411;
	assign w50295 = w15374 ^ w15375;
	assign w50297 = w15402 ^ w15373;
	assign w15486 = w15411 ^ w15385;
	assign w15377 = w15401 ^ w15378;
	assign w15388 = w15392 ^ w44015;
	assign w15387 = w15383 ^ w15388;
	assign w15487 = w15386 ^ w15387;
	assign w15391 = w44019 ^ w15388;
	assign w15488 = w15390 ^ w15391;
	assign w50294 = w15376 ^ w15377;
	assign w45314 = ~w15487;
	assign w45315 = ~w15488;
	assign w45321 = ~w15486;
	assign w29572 = w29667 ^ w29616;
	assign w29654 = w46683 ^ w29572;
	assign w29652 = w29653 & w29654;
	assign w29651 = w29652 ^ w29660;
	assign w29570 = w29652 ^ w29669;
	assign w29628 = w29651 & w29683;
	assign w29571 = w29652 ^ w29616;
	assign w29637 = w29651 & w46684;
	assign w29565 = w29570 ^ w29666;
	assign w29650 = w29658 ^ w29652;
	assign w29649 = w29660 & w29650;
	assign w29647 = w29649 ^ w29657;
	assign w44611 = w29649 ^ w29667;
	assign w29641 = w44611 ^ w29619;
	assign w29639 = w29641 & w29678;
	assign w29630 = w29641 & w29682;
	assign w29608 = w46683 ^ w44611;
	assign w29648 = w29608 ^ w29571;
	assign w29629 = w29648 & w29679;
	assign w29638 = w29648 & w29677;
	assign w44614 = w29637 ^ w29639;
	assign w29643 = w29565 ^ w29566;
	assign w29624 = w29643 & w29686;
	assign w29633 = w29643 & w29675;
	assign w29562 = w46679 ^ w29563;
	assign w29646 = w29655 & w29647;
	assign w29611 = w29646 ^ w29621;
	assign w29569 = w29646 ^ w29670;
	assign w29561 = w29608 ^ w29569;
	assign w29568 = w29598 ^ w29561;
	assign w29640 = w29561 ^ w29562;
	assign w29632 = w29640 & w29673;
	assign w29644 = w29565 ^ w29568;
	assign w29631 = w29644 & w29676;
	assign w29623 = w29640 & w29688;
	assign w29622 = w29644 & w29685;
	assign w29588 = w29633 ^ w29622;
	assign w29584 = ~w29588;
	assign w29645 = w29611 ^ w29613;
	assign w29626 = w29645 & w29680;
	assign w29635 = w29645 & w29684;
	assign w29593 = w29632 ^ w29635;
	assign w29590 = ~w29593;
	assign w29596 = w29634 ^ w29626;
	assign w29578 = w29634 ^ w29635;
	assign w29642 = w29611 ^ w29564;
	assign w29627 = w29642 & w29687;
	assign w29636 = w29642 & w29672;
	assign w29609 = w29627 ^ w29631;
	assign w29587 = ~w29609;
	assign w29594 = w29636 ^ w29627;
	assign w29586 = w29587 ^ w29625;
	assign w29582 = w29586 ^ w44614;
	assign w29585 = w29624 ^ w29582;
	assign w29689 = w29584 ^ w29585;
	assign w44613 = w29635 ^ w29636;
	assign w29617 = w29632 ^ w44613;
	assign w29577 = w29633 ^ w29617;
	assign w29583 = w29628 ^ w29617;
	assign w29580 = ~w29583;
	assign w45681 = ~w29689;
	assign w29589 = w29632 ^ w29633;
	assign w44610 = w29623 ^ w29624;
	assign w29592 = w29596 ^ w44610;
	assign w29591 = w29587 ^ w29592;
	assign w29691 = w29590 ^ w29591;
	assign w45675 = ~w29691;
	assign w29595 = w44614 ^ w29592;
	assign w29692 = w29594 ^ w29595;
	assign w45676 = ~w29692;
	assign w29605 = w29629 ^ w44610;
	assign w29581 = w29605 ^ w29582;
	assign w50279 = w29580 ^ w29581;
	assign w29606 = w29630 ^ w29605;
	assign w50282 = w29606 ^ w29577;
	assign w29610 = w29638 ^ w29606;
	assign w29615 = w29639 ^ w29610;
	assign w50281 = w44613 ^ w29615;
	assign w29579 = w29637 ^ w29610;
	assign w50280 = w29578 ^ w29579;
	assign w29690 = w29615 ^ w29589;
	assign w45674 = ~w29690;
	assign w45941 = ~w9139;
	assign w8971 = w45941 ^ w45610;
	assign w9058 = w45941 ^ w49857;
	assign w49744 = w9057 ^ w9058;
	assign w46840 = w49744 ^ w1082;
	assign w24060 = w46842 ^ w46840;
	assign w24045 = w23970 ^ w24060;
	assign w24058 = w46840 ^ w46837;
	assign w24054 = w24058 ^ w23986;
	assign w8934 = w45941 ^ w49859;
	assign w49723 = w8971 ^ w8972;
	assign w46861 = w49723 ^ w1061;
	assign w27052 = w46863 ^ w46861;
	assign w27127 = w27052 ^ w27142;
	assign w27139 = w46861 ^ w46866;
	assign w27140 = w46864 ^ w46861;
	assign w27136 = w27140 ^ w27068;
	assign w27132 = w27051 ^ w27140;
	assign w27131 = w46868 ^ w27132;
	assign w27125 = w27132 & w27136;
	assign w27057 = w27125 ^ w27054;
	assign w27119 = w27140 & w27129;
	assign w27055 = w27119 ^ w27053;
	assign w27014 = w27054 ^ w27052;
	assign w27130 = w27051 ^ w27014;
	assign w27117 = w27139 & w27130;
	assign w27118 = w27142 & w27127;
	assign w27027 = w27118 ^ w27119;
	assign w27074 = w27027 ^ w27028;
	assign w24036 = w24060 & w24045;
	assign w27135 = w27052 ^ w27058;
	assign w27133 = w27068 ^ w27135;
	assign w27124 = w27133 & w27131;
	assign w27120 = w27135 & w27128;
	assign w44502 = w27117 ^ w27120;
	assign w23972 = w46840 ^ w46838;
	assign w23932 = w23972 ^ w23970;
	assign w23931 = w23972 ^ w46839;
	assign w24055 = w46844 ^ w23931;
	assign w27141 = w46861 ^ w46867;
	assign w27122 = w27141 & w27126;
	assign w27056 = w27122 ^ w27052;
	assign w27073 = w27074 ^ w27056;
	assign w27115 = w27121 ^ w27073;
	assign w27030 = w27056 ^ w44502;
	assign w27114 = w27030 ^ w27055;
	assign w27061 = w27057 ^ w27055;
	assign w27066 = w46861 ^ w27061;
	assign w9207 = w8934 ^ w8935;
	assign w49743 = w9207 ^ w9204;
	assign w46841 = w49743 ^ w1081;
	assign w23969 = w46843 ^ w46841;
	assign w24048 = w23969 ^ w23932;
	assign w24050 = w23969 ^ w24058;
	assign w24043 = w24050 & w24054;
	assign w23975 = w24043 ^ w23972;
	assign w23946 = w46841 ^ w46842;
	assign w24049 = w46844 ^ w24050;
	assign w24042 = w24051 & w24049;
	assign w23993 = w24036 ^ w24042;
	assign w24035 = w24057 & w24048;
	assign w23971 = w46842 ^ w23969;
	assign w24046 = w23976 ^ w23971;
	assign w24044 = w46839 ^ w23971;
	assign w24040 = w24059 & w24044;
	assign w23974 = w24040 ^ w23970;
	assign w24047 = w46838 ^ w23971;
	assign w24038 = w24053 & w24046;
	assign w24037 = w24058 & w24047;
	assign w23973 = w24037 ^ w23971;
	assign w23979 = w23975 ^ w23973;
	assign w23984 = w46837 ^ w23979;
	assign w23945 = w24036 ^ w24037;
	assign w23992 = w23945 ^ w23946;
	assign w23991 = w23992 ^ w23974;
	assign w24033 = w24039 ^ w23991;
	assign w44374 = w24035 ^ w24038;
	assign w23948 = w23974 ^ w44374;
	assign w24032 = w23948 ^ w23973;
	assign w23988 = w24036 ^ w44374;
	assign w23944 = w24039 ^ w23988;
	assign w24026 = w46843 ^ w23944;
	assign w24034 = w23993 ^ w23984;
	assign w24030 = w24034 & w24033;
	assign w24029 = w24030 ^ w24032;
	assign w27070 = w27118 ^ w44502;
	assign w27026 = w27121 ^ w27070;
	assign w27108 = w46867 ^ w27026;
	assign w27075 = w27118 ^ w27124;
	assign w27116 = w27075 ^ w27066;
	assign w27112 = w27116 & w27115;
	assign w27111 = w27112 ^ w27114;
	assign w44501 = w27117 ^ w27123;
	assign w27029 = w27061 ^ w44501;
	assign w27072 = w46863 ^ w27029;
	assign w27107 = w27112 ^ w27072;
	assign w27106 = w27107 & w27108;
	assign w27104 = w27112 ^ w27106;
	assign w27025 = w27106 ^ w27070;
	assign w27024 = w27106 ^ w27123;
	assign w27019 = w27024 ^ w27120;
	assign w27103 = w27114 & w27104;
	assign w27101 = w27103 ^ w27111;
	assign w44505 = w27103 ^ w27121;
	assign w27095 = w44505 ^ w27073;
	assign w27084 = w27095 & w27136;
	assign w27093 = w27095 & w27132;
	assign w27062 = w46867 ^ w44505;
	assign w27102 = w27062 ^ w27025;
	assign w27083 = w27102 & w27133;
	assign w27092 = w27102 & w27131;
	assign w27105 = w27106 ^ w27114;
	assign w27091 = w27105 & w46868;
	assign w27082 = w27105 & w27137;
	assign w44504 = w27091 ^ w27093;
	assign w27067 = w44501 ^ w27052;
	assign w27113 = w27075 ^ w27067;
	assign w27110 = w27113 & w27111;
	assign w27018 = w27110 ^ w27066;
	assign w27109 = w27110 ^ w27072;
	assign w27088 = w27109 & w27128;
	assign w27079 = w27109 & w27135;
	assign w27021 = w27110 ^ w27122;
	assign w27017 = w27021 ^ w27057;
	assign w27016 = w46863 ^ w27017;
	assign w27020 = w46861 ^ w27017;
	assign w27097 = w27019 ^ w27020;
	assign w27078 = w27097 & w27140;
	assign w27087 = w27097 & w27129;
	assign w24041 = w46844 & w24055;
	assign w44377 = w24035 ^ w24041;
	assign w23947 = w23979 ^ w44377;
	assign w23990 = w46839 ^ w23947;
	assign w24025 = w24030 ^ w23990;
	assign w24024 = w24025 & w24026;
	assign w24022 = w24030 ^ w24024;
	assign w24021 = w24032 & w24022;
	assign w24019 = w24021 ^ w24029;
	assign w24023 = w24024 ^ w24032;
	assign w24009 = w24023 & w46844;
	assign w24000 = w24023 & w24055;
	assign w23942 = w24024 ^ w24041;
	assign w23937 = w23942 ^ w24038;
	assign w44376 = w24021 ^ w24039;
	assign w23980 = w46843 ^ w44376;
	assign w24013 = w44376 ^ w23991;
	assign w24011 = w24013 & w24050;
	assign w24002 = w24013 & w24054;
	assign w44379 = w24009 ^ w24011;
	assign w23985 = w44377 ^ w23970;
	assign w24031 = w23993 ^ w23985;
	assign w24028 = w24031 & w24029;
	assign w23936 = w24028 ^ w23984;
	assign w24027 = w24028 ^ w23990;
	assign w23997 = w24027 & w24053;
	assign w23939 = w24028 ^ w24040;
	assign w23935 = w23939 ^ w23975;
	assign w23938 = w46837 ^ w23935;
	assign w24015 = w23937 ^ w23938;
	assign w23996 = w24015 & w24058;
	assign w24005 = w24015 & w24047;
	assign w24018 = w24027 & w24019;
	assign w23941 = w24018 ^ w24042;
	assign w23933 = w23980 ^ w23941;
	assign w23983 = w24018 ^ w23993;
	assign w24017 = w23983 ^ w23985;
	assign w23998 = w24017 & w24052;
	assign w24007 = w24017 & w24056;
	assign w24006 = w24027 & w24046;
	assign w23968 = w24006 ^ w23998;
	assign w23950 = w24006 ^ w24007;
	assign w23934 = w46839 ^ w23935;
	assign w24012 = w23933 ^ w23934;
	assign w24004 = w24012 & w24045;
	assign w23961 = w24004 ^ w24005;
	assign w23965 = w24004 ^ w24007;
	assign w23962 = ~w23965;
	assign w23995 = w24012 & w24060;
	assign w44375 = w23995 ^ w23996;
	assign w23964 = w23968 ^ w44375;
	assign w23967 = w44379 ^ w23964;
	assign w23940 = w23970 ^ w23933;
	assign w24016 = w23937 ^ w23940;
	assign w23994 = w24016 & w24057;
	assign w24003 = w24016 & w24048;
	assign w23960 = w24005 ^ w23994;
	assign w23956 = ~w23960;
	assign w23943 = w24024 ^ w23988;
	assign w24020 = w23980 ^ w23943;
	assign w24001 = w24020 & w24051;
	assign w23977 = w24001 ^ w44375;
	assign w23978 = w24002 ^ w23977;
	assign w24010 = w24020 & w24049;
	assign w23982 = w24010 ^ w23978;
	assign w23951 = w24009 ^ w23982;
	assign w23987 = w24011 ^ w23982;
	assign w24062 = w23987 ^ w23961;
	assign w50063 = ~w24062;
	assign w9529 = w45327 ^ w50063;
	assign w9336 = w9529 ^ w45338;
	assign w9398 = w9529 ^ w9485;
	assign w49948 = w50059 ^ w9398;
	assign w9411 = w9535 ^ w24062;
	assign w9427 = w9537 ^ w9529;
	assign w49931 = w45339 ^ w9427;
	assign w49939 = w9411 ^ w9412;
	assign w46709 = w49948 ^ w1213;
	assign w46718 = w49939 ^ w1204;
	assign w46726 = w49931 ^ w1196;
	assign w50061 = w23950 ^ w23951;
	assign w9235 = w50061 ^ w50051;
	assign w9539 = w50057 ^ w50061;
	assign w9419 = w9420 ^ w50061;
	assign w49936 = w9418 ^ w9419;
	assign w46721 = w49936 ^ w1201;
	assign w9317 = w24062 ^ w50054;
	assign w9404 = w9540 ^ w9539;
	assign w9402 = ~w9404;
	assign w49928 = w9554 ^ w9539;
	assign w46729 = w49928 ^ w1193;
	assign w27100 = w27109 & w27101;
	assign w27023 = w27100 ^ w27124;
	assign w27015 = w27062 ^ w27023;
	assign w27022 = w27052 ^ w27015;
	assign w27098 = w27019 ^ w27022;
	assign w27076 = w27098 & w27139;
	assign w27094 = w27015 ^ w27016;
	assign w27077 = w27094 & w27142;
	assign w27086 = w27094 & w27127;
	assign w27085 = w27098 & w27130;
	assign w27043 = w27086 ^ w27087;
	assign w43576 = w27077 ^ w27078;
	assign w27059 = w27083 ^ w43576;
	assign w27060 = w27084 ^ w27059;
	assign w27064 = w27092 ^ w27060;
	assign w27069 = w27093 ^ w27064;
	assign w27144 = w27069 ^ w27043;
	assign w50104 = ~w27144;
	assign w27042 = w27087 ^ w27076;
	assign w27038 = ~w27042;
	assign w27065 = w27100 ^ w27075;
	assign w27096 = w27065 ^ w27018;
	assign w27081 = w27096 & w27141;
	assign w27063 = w27081 ^ w27085;
	assign w27041 = ~w27063;
	assign w27090 = w27096 & w27126;
	assign w27048 = w27090 ^ w27081;
	assign w27099 = w27065 ^ w27067;
	assign w27080 = w27099 & w27134;
	assign w27050 = w27088 ^ w27080;
	assign w27046 = w27050 ^ w43576;
	assign w27045 = w27041 ^ w27046;
	assign w27049 = w44504 ^ w27046;
	assign w27146 = w27048 ^ w27049;
	assign w27040 = w27041 ^ w27079;
	assign w27036 = w27040 ^ w44504;
	assign w27035 = w27059 ^ w27036;
	assign w27039 = w27078 ^ w27036;
	assign w27143 = w27038 ^ w27039;
	assign w27089 = w27099 & w27138;
	assign w27032 = w27088 ^ w27089;
	assign w27047 = w27086 ^ w27089;
	assign w27044 = ~w27047;
	assign w27145 = w27044 ^ w27045;
	assign w44503 = w27089 ^ w27090;
	assign w27071 = w27086 ^ w44503;
	assign w27037 = w27082 ^ w27071;
	assign w27031 = w27087 ^ w27071;
	assign w50105 = w27060 ^ w27031;
	assign w9490 = w50105 ^ w50117;
	assign w9289 = w9528 ^ w9490;
	assign w50103 = w44503 ^ w27069;
	assign w9284 = ~w50103;
	assign w9473 = w50116 ^ w9284;
	assign w45602 = ~w27145;
	assign w9287 = w9496 ^ w45602;
	assign w45603 = ~w27146;
	assign w9244 = w9490 ^ w45603;
	assign w45609 = ~w27143;
	assign w9457 = w27144 ^ w45609;
	assign w9513 = w45609 ^ w45521;
	assign w9447 = w9513 ^ w50112;
	assign w9471 = w9513 ^ w9501;
	assign w27034 = ~w27037;
	assign w50101 = w27034 ^ w27035;
	assign w9246 = w9490 ^ w50101;
	assign w9566 = w9246 ^ w9247;
	assign w27033 = w27091 ^ w27064;
	assign w50102 = w27032 ^ w27033;
	assign w9504 = w50102 ^ w50115;
	assign w9475 = w9504 ^ w9495;
	assign w24014 = w23983 ^ w23936;
	assign w23999 = w24014 & w24059;
	assign w24008 = w24014 & w24044;
	assign w23981 = w23999 ^ w24003;
	assign w44378 = w24007 ^ w24008;
	assign w50062 = w44378 ^ w23987;
	assign w9536 = w50058 ^ w50062;
	assign w9401 = w9537 ^ w9536;
	assign w49946 = w45326 ^ w9401;
	assign w46711 = w49946 ^ w1211;
	assign w29732 = w46711 ^ w46709;
	assign w9429 = w9431 ^ w9536;
	assign w23989 = w24004 ^ w44378;
	assign w23949 = w24005 ^ w23989;
	assign w50064 = w23978 ^ w23949;
	assign w9492 = w50048 ^ w50064;
	assign w9234 = w9492 ^ w50046;
	assign w9571 = w9234 ^ w9235;
	assign w9477 = w9525 ^ w9492;
	assign w9388 = ~w9492;
	assign w9387 = w9388 ^ w50050;
	assign w49921 = w9571 ^ w9536;
	assign w46736 = w49921 ^ w1186;
	assign w9484 = w50059 ^ w50064;
	assign w9426 = w9535 ^ w9484;
	assign w49932 = w50048 ^ w9426;
	assign w46725 = w49932 ^ w1197;
	assign w9408 = w9525 ^ w9484;
	assign w49941 = w45341 ^ w9408;
	assign w46716 = w49941 ^ w1206;
	assign w23959 = ~w23981;
	assign w23963 = w23959 ^ w23964;
	assign w23958 = w23959 ^ w23997;
	assign w24063 = w23962 ^ w23963;
	assign w23954 = w23958 ^ w44379;
	assign w23957 = w23996 ^ w23954;
	assign w24061 = w23956 ^ w23957;
	assign w23966 = w24008 ^ w23999;
	assign w24064 = w23966 ^ w23967;
	assign w9354 = w50062 ^ w33173;
	assign w9271 = w9486 ^ w50062;
	assign w45518 = ~w24061;
	assign w9532 = w45326 ^ w45518;
	assign w9355 = w9532 ^ w50047;
	assign w9353 = ~w9355;
	assign w49922 = w9353 ^ w9354;
	assign w9399 = w9535 ^ w9532;
	assign w49947 = w45327 ^ w9399;
	assign w9413 = w9537 ^ w45518;
	assign w49938 = w9413 ^ w9414;
	assign w9428 = w9540 ^ w9532;
	assign w49930 = w45338 ^ w9428;
	assign w46735 = w49922 ^ w1187;
	assign w46719 = w49938 ^ w1203;
	assign w46710 = w49947 ^ w1212;
	assign w9337 = w45518 ^ w33174;
	assign w9335 = w9336 ^ w9337;
	assign w49923 = ~w9335;
	assign w46734 = w49923 ^ w1188;
	assign w29738 = w46716 ^ w46710;
	assign w29818 = w46711 ^ w29738;
	assign w29815 = w29732 ^ w29738;
	assign w46727 = w49930 ^ w1195;
	assign w11374 = w46727 ^ w46725;
	assign w45519 = ~w24063;
	assign w9417 = w9388 ^ w45519;
	assign w9406 = w45519 ^ w15889;
	assign w49943 = w9405 ^ w9406;
	assign w46714 = w49943 ^ w1208;
	assign w29819 = w46709 ^ w46714;
	assign w9547 = w45340 ^ w45519;
	assign w9423 = w9547 ^ w9525;
	assign w9422 = w9423 ^ w9424;
	assign w49934 = ~w9422;
	assign w9400 = w9547 ^ w9524;
	assign w46723 = w49934 ^ w1199;
	assign w26649 = w46723 ^ w46721;
	assign w45520 = ~w24064;
	assign w9277 = w9484 ^ w45520;
	assign w9553 = w9277 ^ w9278;
	assign w49917 = w45520 ^ w9477;
	assign w46740 = w49917 ^ w1182;
	assign w15668 = w46740 ^ w46734;
	assign w15748 = w46735 ^ w15668;
	assign w9548 = w45341 ^ w45520;
	assign w9416 = w9548 ^ w9526;
	assign w9415 = w9416 ^ w9417;
	assign w9425 = w9548 ^ w9486;
	assign w49918 = ~w9415;
	assign w49933 = w45766 ^ w9425;
	assign w9300 = w9548 ^ w9485;
	assign w46739 = w49918 ^ w1183;
	assign w15744 = w46739 ^ w15748;
	assign w15731 = w15748 & w15744;
	assign w46724 = w49933 ^ w1198;
	assign w49925 = w45328 ^ w9300;
	assign w46732 = w49925 ^ w1190;
	assign w11380 = w46732 ^ w46726;
	assign w11457 = w11374 ^ w11380;
	assign w49942 = w9553 ^ w9526;
	assign w46715 = w49942 ^ w1207;
	assign w29748 = w46715 ^ w46714;
	assign w29813 = w29748 ^ w29815;
	assign w29821 = w46709 ^ w46715;
	assign w29814 = w46715 ^ w29818;
	assign w29801 = w29818 & w29814;
	assign w26656 = w46724 ^ w46718;
	assign w26736 = w46719 ^ w26656;
	assign w26732 = w46723 ^ w26736;
	assign w26719 = w26736 & w26732;
	assign w9556 = w9271 ^ w9272;
	assign w49937 = w9556 ^ w9540;
	assign w46720 = w49937 ^ w1202;
	assign w26652 = w46720 ^ w46718;
	assign w26611 = w26652 ^ w46719;
	assign w26735 = w46724 ^ w26611;
	assign w26721 = w46724 & w26735;
	assign w11460 = w46727 ^ w11380;
	assign w23955 = w24000 ^ w23989;
	assign w23952 = ~w23955;
	assign w15664 = w46736 ^ w46734;
	assign w15623 = w15664 ^ w46735;
	assign w15747 = w46740 ^ w15623;
	assign w15733 = w46740 & w15747;
	assign w23953 = w23977 ^ w23954;
	assign w50060 = w23952 ^ w23953;
	assign w9527 = w50045 ^ w50060;
	assign w49919 = w50060 ^ w9400;
	assign w9421 = w9527 ^ w9526;
	assign w49935 = w50049 ^ w9421;
	assign w9389 = ~w9527;
	assign w46722 = w49935 ^ w1200;
	assign w26666 = w46723 ^ w46722;
	assign w26740 = w46722 ^ w46720;
	assign w26651 = w46722 ^ w26649;
	assign w26727 = w46718 ^ w26651;
	assign w26724 = w46719 ^ w26651;
	assign w9386 = w9539 ^ w9389;
	assign w49920 = w9386 ^ w9387;
	assign w46737 = w49920 ^ w1185;
	assign w15661 = w46739 ^ w46737;
	assign w26626 = w46721 ^ w46722;
	assign w9458 = w9389 ^ w45773;
	assign w49927 = w9458 ^ w9459;
	assign w46730 = w49927 ^ w1192;
	assign w11350 = w46729 ^ w46730;
	assign w46738 = w49919 ^ w1184;
	assign w15663 = w46738 ^ w15661;
	assign w15736 = w46735 ^ w15663;
	assign w15738 = w15668 ^ w15663;
	assign w15739 = w46734 ^ w15663;
	assign w15678 = w46739 ^ w46738;
	assign w15752 = w46738 ^ w46736;
	assign w26726 = w26656 ^ w26651;
	assign w15638 = w46737 ^ w46738;
	assign w11461 = w46725 ^ w46730;
	assign w45942 = ~w9137;
	assign w9035 = w45942 ^ w49865;
	assign w9039 = w45942 ^ w45357;
	assign w49759 = w9034 ^ w9035;
	assign w46825 = w49759 ^ w1033;
	assign w11618 = w46825 ^ w46826;
	assign w9037 = w9038 ^ w9039;
	assign w49757 = ~w9037;
	assign w46827 = w49757 ^ w1031;
	assign w11641 = w46827 ^ w46825;
	assign w11724 = w46827 ^ w11728;
	assign w11711 = w11728 & w11724;
	assign w9032 = w45942 ^ w49866;
	assign w49760 = w9031 ^ w9032;
	assign w46824 = w49760 ^ w1034;
	assign w11732 = w46826 ^ w46824;
	assign w11644 = w46824 ^ w46822;
	assign w11604 = w11644 ^ w11642;
	assign w11603 = w11644 ^ w46823;
	assign w11730 = w46824 ^ w46821;
	assign w11658 = w46827 ^ w46826;
	assign w11726 = w11730 ^ w11658;
	assign w11722 = w11641 ^ w11730;
	assign w11721 = w46828 ^ w11722;
	assign w11731 = w46821 ^ w46827;
	assign w11715 = w11722 & w11726;
	assign w11647 = w11715 ^ w11644;
	assign w11717 = w11642 ^ w11732;
	assign w11708 = w11732 & w11717;
	assign w11723 = w11658 ^ w11725;
	assign w11714 = w11723 & w11721;
	assign w11665 = w11708 ^ w11714;
	assign w11643 = w46826 ^ w11641;
	assign w11719 = w46822 ^ w11643;
	assign w11716 = w46823 ^ w11643;
	assign w11712 = w11731 & w11716;
	assign w11709 = w11730 & w11719;
	assign w11718 = w11648 ^ w11643;
	assign w11710 = w11725 & w11718;
	assign w11645 = w11709 ^ w11643;
	assign w11617 = w11708 ^ w11709;
	assign w11664 = w11617 ^ w11618;
	assign w11651 = w11647 ^ w11645;
	assign w11646 = w11712 ^ w11642;
	assign w11663 = w11664 ^ w11646;
	assign w11705 = w11711 ^ w11663;
	assign w11656 = w46821 ^ w11651;
	assign w11706 = w11665 ^ w11656;
	assign w11702 = w11706 & w11705;
	assign w11720 = w11641 ^ w11604;
	assign w11707 = w11729 & w11720;
	assign w43858 = w11707 ^ w11710;
	assign w11660 = w11708 ^ w43858;
	assign w11616 = w11711 ^ w11660;
	assign w11698 = w46827 ^ w11616;
	assign w11727 = w46828 ^ w11603;
	assign w11713 = w46828 & w11727;
	assign w43861 = w11707 ^ w11713;
	assign w11619 = w11651 ^ w43861;
	assign w11662 = w46823 ^ w11619;
	assign w11697 = w11702 ^ w11662;
	assign w11696 = w11697 & w11698;
	assign w11694 = w11702 ^ w11696;
	assign w11614 = w11696 ^ w11713;
	assign w11609 = w11614 ^ w11710;
	assign w11657 = w43861 ^ w11642;
	assign w11703 = w11665 ^ w11657;
	assign w11615 = w11696 ^ w11660;
	assign w11620 = w11646 ^ w43858;
	assign w11704 = w11620 ^ w11645;
	assign w11695 = w11696 ^ w11704;
	assign w11681 = w11695 & w46828;
	assign w11672 = w11695 & w11727;
	assign w11693 = w11704 & w11694;
	assign w43860 = w11693 ^ w11711;
	assign w11685 = w43860 ^ w11663;
	assign w11674 = w11685 & w11726;
	assign w11683 = w11685 & w11722;
	assign w43863 = w11681 ^ w11683;
	assign w11701 = w11702 ^ w11704;
	assign w11700 = w11703 & w11701;
	assign w11691 = w11693 ^ w11701;
	assign w11611 = w11700 ^ w11712;
	assign w11607 = w11611 ^ w11647;
	assign w11606 = w46823 ^ w11607;
	assign w11652 = w46827 ^ w43860;
	assign w11692 = w11652 ^ w11615;
	assign w11682 = w11692 & w11721;
	assign w11673 = w11692 & w11723;
	assign w11699 = w11700 ^ w11662;
	assign w11669 = w11699 & w11725;
	assign w11678 = w11699 & w11718;
	assign w11690 = w11699 & w11691;
	assign w11613 = w11690 ^ w11714;
	assign w11655 = w11690 ^ w11665;
	assign w11689 = w11655 ^ w11657;
	assign w11679 = w11689 & w11728;
	assign w11622 = w11678 ^ w11679;
	assign w11670 = w11689 & w11724;
	assign w11640 = w11678 ^ w11670;
	assign w11605 = w11652 ^ w11613;
	assign w11612 = w11642 ^ w11605;
	assign w11688 = w11609 ^ w11612;
	assign w11666 = w11688 & w11729;
	assign w11675 = w11688 & w11720;
	assign w11684 = w11605 ^ w11606;
	assign w11667 = w11684 & w11732;
	assign w11676 = w11684 & w11717;
	assign w11637 = w11676 ^ w11679;
	assign w11634 = ~w11637;
	assign w11610 = w46821 ^ w11607;
	assign w11687 = w11609 ^ w11610;
	assign w11668 = w11687 & w11730;
	assign w11677 = w11687 & w11719;
	assign w11632 = w11677 ^ w11666;
	assign w11628 = ~w11632;
	assign w43859 = w11667 ^ w11668;
	assign w11636 = w11640 ^ w43859;
	assign w11639 = w43863 ^ w11636;
	assign w11633 = w11676 ^ w11677;
	assign w11649 = w11673 ^ w43859;
	assign w11650 = w11674 ^ w11649;
	assign w11654 = w11682 ^ w11650;
	assign w11623 = w11681 ^ w11654;
	assign w50107 = w11622 ^ w11623;
	assign w9283 = w50107 ^ w9284;
	assign w11659 = w11683 ^ w11654;
	assign w9498 = w50107 ^ w50111;
	assign w9437 = w9498 ^ w9496;
	assign w50016 = w9566 ^ w9498;
	assign w46641 = w50016 ^ w1089;
	assign w11734 = w11659 ^ w11633;
	assign w45236 = ~w11734;
	assign w50019 = w45236 ^ w9471;
	assign w9543 = w50104 ^ w45236;
	assign w9445 = w45331 ^ w45236;
	assign w9454 = w9543 ^ w9478;
	assign w50028 = w50105 ^ w9454;
	assign w9433 = w9543 ^ w45521;
	assign w46629 = w50028 ^ w1101;
	assign w46638 = w50019 ^ w1092;
	assign w50043 = w9433 ^ w9434;
	assign w46614 = w50043 ^ w1116;
	assign w11608 = w11700 ^ w11656;
	assign w11686 = w11655 ^ w11608;
	assign w11680 = w11686 & w11716;
	assign w11671 = w11686 & w11731;
	assign w11653 = w11671 ^ w11675;
	assign w11638 = w11680 ^ w11671;
	assign w43862 = w11679 ^ w11680;
	assign w50108 = w43862 ^ w11659;
	assign w9544 = w50103 ^ w50108;
	assign w9460 = w9544 ^ w9513;
	assign w50026 = w45330 ^ w9460;
	assign w9449 = w9544 ^ w9498;
	assign w46631 = w50026 ^ w1099;
	assign w11106 = w46631 ^ w46629;
	assign w50041 = w9550 ^ w9544;
	assign w46616 = w50041 ^ w1114;
	assign w29466 = w46616 ^ w46614;
	assign w9476 = w9490 ^ w50108;
	assign w50017 = w9475 ^ w9476;
	assign w46640 = w50017 ^ w1090;
	assign w15128 = w46640 ^ w46638;
	assign w11661 = w11676 ^ w43862;
	assign w11621 = w11677 ^ w11661;
	assign w11627 = w11672 ^ w11661;
	assign w11624 = ~w11627;
	assign w50109 = w11650 ^ w11621;
	assign w9493 = w50109 ^ w50113;
	assign w9232 = w9493 ^ w50110;
	assign w9230 = w9493 ^ w45515;
	assign w9470 = w50109 ^ w27144;
	assign w9450 = w9493 ^ w50116;
	assign w50033 = w9449 ^ w9450;
	assign w46624 = w50033 ^ w1106;
	assign w9479 = w50105 ^ w50109;
	assign w9468 = w9528 ^ w9479;
	assign w9444 = w9479 ^ w50117;
	assign w50021 = w45603 ^ w9468;
	assign w50036 = w9444 ^ w9445;
	assign w46621 = w50036 ^ w1109;
	assign w26470 = w46624 ^ w46621;
	assign w46636 = w50021 ^ w1094;
	assign w11631 = ~w11653;
	assign w11630 = w11631 ^ w11669;
	assign w11626 = w11630 ^ w43863;
	assign w11629 = w11668 ^ w11626;
	assign w11733 = w11628 ^ w11629;
	assign w11625 = w11649 ^ w11626;
	assign w50106 = w11624 ^ w11625;
	assign w9233 = w50107 ^ w50106;
	assign w9572 = w9232 ^ w9233;
	assign w9288 = w45515 ^ w50106;
	assign w50015 = w9287 ^ w9288;
	assign w46642 = w50015 ^ w1088;
	assign w15102 = w46641 ^ w46642;
	assign w50032 = w9572 ^ w9504;
	assign w46625 = w50032 ^ w1105;
	assign w9518 = w50101 ^ w50106;
	assign w9439 = w9518 ^ w9508;
	assign w9451 = w9518 ^ w50114;
	assign w9463 = w9518 ^ w9504;
	assign w9461 = ~w9463;
	assign w50039 = w50110 ^ w9439;
	assign w46618 = w50039 ^ w1112;
	assign w29554 = w46618 ^ w46616;
	assign w9432 = w9501 ^ w9479;
	assign w50044 = w50113 ^ w9432;
	assign w46613 = w50044 ^ w1117;
	assign w29552 = w46616 ^ w46613;
	assign w15216 = w46642 ^ w46640;
	assign w11736 = w11638 ^ w11639;
	assign w45230 = ~w11736;
	assign w9541 = w45603 ^ w45230;
	assign w9466 = w9541 ^ w9508;
	assign w9453 = w9541 ^ w9493;
	assign w50029 = w45516 ^ w9453;
	assign w9443 = w9541 ^ w9478;
	assign w50037 = w45333 ^ w9443;
	assign w50013 = w45230 ^ w9289;
	assign w9231 = w45333 ^ w45230;
	assign w9573 = w9230 ^ w9231;
	assign w46644 = w50013 ^ w1086;
	assign w15132 = w46644 ^ w46638;
	assign w46620 = w50037 ^ w1110;
	assign w29470 = w46620 ^ w46614;
	assign w46628 = w50029 ^ w1102;
	assign w45235 = ~w11733;
	assign w9448 = w45235 ^ w50108;
	assign w9456 = w9501 ^ w45235;
	assign w9455 = w9456 ^ w9457;
	assign w50027 = ~w9455;
	assign w50034 = w9447 ^ w9448;
	assign w46623 = w50034 ^ w1107;
	assign w9503 = w45235 ^ w45330;
	assign w9474 = ~w9503;
	assign w9446 = w9543 ^ w9503;
	assign w50035 = w45514 ^ w9446;
	assign w9472 = w9474 ^ w45521;
	assign w50018 = w9472 ^ w9473;
	assign w9435 = w9503 ^ w9495;
	assign w50042 = w45609 ^ w9435;
	assign w26382 = w46623 ^ w46621;
	assign w46639 = w50018 ^ w1091;
	assign w15212 = w46639 ^ w15132;
	assign w46622 = w50035 ^ w1108;
	assign w26388 = w46628 ^ w46622;
	assign w26468 = w46623 ^ w26388;
	assign w26384 = w46624 ^ w46622;
	assign w26344 = w26384 ^ w26382;
	assign w26343 = w26384 ^ w46623;
	assign w26467 = w46628 ^ w26343;
	assign w26453 = w46628 & w26467;
	assign w46630 = w50027 ^ w1100;
	assign w46615 = w50042 ^ w1115;
	assign w29550 = w46615 ^ w29470;
	assign w26465 = w26382 ^ w26388;
	assign w11112 = w46636 ^ w46630;
	assign w11192 = w46631 ^ w11112;
	assign w11189 = w11106 ^ w11112;
	assign w29464 = w46615 ^ w46613;
	assign w29547 = w29464 ^ w29470;
	assign w29539 = w29464 ^ w29554;
	assign w29530 = w29554 & w29539;
	assign w29426 = w29466 ^ w29464;
	assign w15087 = w15128 ^ w46639;
	assign w15211 = w46644 ^ w15087;
	assign w15197 = w46644 & w15211;
	assign w29425 = w29466 ^ w46615;
	assign w29549 = w46620 ^ w29425;
	assign w29551 = w46613 ^ w46618;
	assign w11635 = w11631 ^ w11636;
	assign w11735 = w11634 ^ w11635;
	assign w45237 = ~w11735;
	assign w9245 = w45516 ^ w45237;
	assign w9452 = w45332 ^ w45237;
	assign w50031 = w9451 ^ w9452;
	assign w9533 = w45602 ^ w45237;
	assign w9464 = w9533 ^ w9496;
	assign w50023 = w50101 ^ w9464;
	assign w9442 = ~w9533;
	assign w9440 = w9442 ^ w9528;
	assign w46626 = w50031 ^ w1104;
	assign w26469 = w46621 ^ w46626;
	assign w26472 = w46626 ^ w46624;
	assign w26358 = w46625 ^ w46626;
	assign w26457 = w26382 ^ w26472;
	assign w26448 = w26472 & w26457;
	assign w46634 = w50023 ^ w1096;
	assign w50030 = w9573 ^ w9533;
	assign w46627 = w50030 ^ w1103;
	assign w26471 = w46621 ^ w46627;
	assign w26398 = w46627 ^ w46626;
	assign w26463 = w26398 ^ w26465;
	assign w26464 = w46627 ^ w26468;
	assign w26451 = w26468 & w26464;
	assign w26466 = w26470 ^ w26398;
	assign w26381 = w46627 ^ w46625;
	assign w26383 = w46626 ^ w26381;
	assign w26460 = w26381 ^ w26344;
	assign w26447 = w26469 & w26460;
	assign w26462 = w26381 ^ w26470;
	assign w26455 = w26462 & w26466;
	assign w26387 = w26455 ^ w26384;
	assign w26461 = w46628 ^ w26462;
	assign w26454 = w26463 & w26461;
	assign w26456 = w46623 ^ w26383;
	assign w26405 = w26448 ^ w26454;
	assign w26459 = w46622 ^ w26383;
	assign w26449 = w26470 & w26459;
	assign w26357 = w26448 ^ w26449;
	assign w26404 = w26357 ^ w26358;
	assign w26385 = w26449 ^ w26383;
	assign w26391 = w26387 ^ w26385;
	assign w26396 = w46621 ^ w26391;
	assign w26446 = w26405 ^ w26396;
	assign w26458 = w26388 ^ w26383;
	assign w26450 = w26465 & w26458;
	assign w44474 = w26447 ^ w26453;
	assign w26397 = w44474 ^ w26382;
	assign w26443 = w26405 ^ w26397;
	assign w26359 = w26391 ^ w44474;
	assign w26402 = w46623 ^ w26359;
	assign w44475 = w26447 ^ w26450;
	assign w26400 = w26448 ^ w44475;
	assign w26356 = w26451 ^ w26400;
	assign w26438 = w46627 ^ w26356;
	assign w9567 = w9244 ^ w9245;
	assign w50014 = w9567 ^ w9508;
	assign w46643 = w50014 ^ w1087;
	assign w15208 = w46643 ^ w15212;
	assign w15142 = w46643 ^ w46642;
	assign w15125 = w46643 ^ w46641;
	assign w15127 = w46642 ^ w15125;
	assign w15203 = w46638 ^ w15127;
	assign w15200 = w46639 ^ w15127;
	assign w15202 = w15132 ^ w15127;
	assign w26452 = w26471 & w26456;
	assign w26386 = w26452 ^ w26382;
	assign w26360 = w26386 ^ w44475;
	assign w26444 = w26360 ^ w26385;
	assign w26403 = w26404 ^ w26386;
	assign w26445 = w26451 ^ w26403;
	assign w26442 = w26446 & w26445;
	assign w26441 = w26442 ^ w26444;
	assign w26440 = w26443 & w26441;
	assign w26437 = w26442 ^ w26402;
	assign w26436 = w26437 & w26438;
	assign w26435 = w26436 ^ w26444;
	assign w26354 = w26436 ^ w26453;
	assign w26412 = w26435 & w26467;
	assign w26355 = w26436 ^ w26400;
	assign w26348 = w26440 ^ w26396;
	assign w26421 = w26435 & w46628;
	assign w26434 = w26442 ^ w26436;
	assign w26433 = w26444 & w26434;
	assign w26431 = w26433 ^ w26441;
	assign w26349 = w26354 ^ w26450;
	assign w26351 = w26440 ^ w26452;
	assign w44478 = w26433 ^ w26451;
	assign w26392 = w46627 ^ w44478;
	assign w26432 = w26392 ^ w26355;
	assign w26413 = w26432 & w26463;
	assign w26425 = w44478 ^ w26403;
	assign w26423 = w26425 & w26462;
	assign w26414 = w26425 & w26466;
	assign w44477 = w26421 ^ w26423;
	assign w26347 = w26351 ^ w26387;
	assign w26350 = w46621 ^ w26347;
	assign w26346 = w46623 ^ w26347;
	assign w26427 = w26349 ^ w26350;
	assign w26408 = w26427 & w26470;
	assign w26417 = w26427 & w26459;
	assign w26439 = w26440 ^ w26402;
	assign w26409 = w26439 & w26465;
	assign w26430 = w26439 & w26431;
	assign w26395 = w26430 ^ w26405;
	assign w26426 = w26395 ^ w26348;
	assign w26429 = w26395 ^ w26397;
	assign w26420 = w26426 & w26456;
	assign w26411 = w26426 & w26471;
	assign w26410 = w26429 & w26464;
	assign w26378 = w26420 ^ w26411;
	assign w26419 = w26429 & w26468;
	assign w26418 = w26439 & w26458;
	assign w26362 = w26418 ^ w26419;
	assign w26380 = w26418 ^ w26410;
	assign w26353 = w26430 ^ w26454;
	assign w26345 = w26392 ^ w26353;
	assign w26424 = w26345 ^ w26346;
	assign w26407 = w26424 & w26472;
	assign w26416 = w26424 & w26457;
	assign w26373 = w26416 ^ w26417;
	assign w26377 = w26416 ^ w26419;
	assign w26374 = ~w26377;
	assign w43573 = w26407 ^ w26408;
	assign w26389 = w26413 ^ w43573;
	assign w26390 = w26414 ^ w26389;
	assign w26376 = w26380 ^ w43573;
	assign w26379 = w44477 ^ w26376;
	assign w26476 = w26378 ^ w26379;
	assign w26352 = w26382 ^ w26345;
	assign w26428 = w26349 ^ w26352;
	assign w26406 = w26428 & w26469;
	assign w26372 = w26417 ^ w26406;
	assign w26368 = ~w26372;
	assign w26415 = w26428 & w26460;
	assign w26393 = w26411 ^ w26415;
	assign w26371 = ~w26393;
	assign w26370 = w26371 ^ w26409;
	assign w26366 = w26370 ^ w44477;
	assign w26365 = w26389 ^ w26366;
	assign w26369 = w26408 ^ w26366;
	assign w26473 = w26368 ^ w26369;
	assign w26375 = w26371 ^ w26376;
	assign w26475 = w26374 ^ w26375;
	assign w50256 = ~w26475;
	assign w43213 = w26475 ^ w45319;
	assign w44476 = w26419 ^ w26420;
	assign w26401 = w26416 ^ w44476;
	assign w26367 = w26412 ^ w26401;
	assign w26364 = ~w26367;
	assign w50257 = w26364 ^ w26365;
	assign w43220 = ~w50257;
	assign w43398 = w45318 ^ w43220;
	assign w26361 = w26417 ^ w26401;
	assign w50260 = w26390 ^ w26361;
	assign w26422 = w26432 & w26461;
	assign w26394 = w26422 ^ w26390;
	assign w26363 = w26421 ^ w26394;
	assign w50258 = w26362 ^ w26363;
	assign w26399 = w26423 ^ w26394;
	assign w26474 = w26399 ^ w26373;
	assign w50259 = w44476 ^ w26399;
	assign w43219 = w50258 ^ w43220;
	assign w15195 = w15212 & w15208;
	assign w45582 = ~w26476;
	assign w43217 = w45318 ^ w45582;
	assign w45588 = ~w26473;
	assign w45589 = ~w26474;
	assign w11193 = w46629 ^ w46634;
	assign w29535 = w46620 & w29549;
	assign w45943 = ~w9135;
	assign w8949 = w45943 ^ w49894;
	assign w49808 = w8948 ^ w8949;
	assign w46776 = w49808 ^ w1018;
	assign w8957 = w45943 ^ w45361;
	assign w49805 = w8956 ^ w8957;
	assign w46779 = w49805 ^ w1015;
	assign w29882 = w46779 ^ w46778;
	assign w29955 = w46773 ^ w46779;
	assign w29947 = w29882 ^ w29949;
	assign w8952 = w45943 ^ w49893;
	assign w29868 = w46776 ^ w46774;
	assign w29827 = w29868 ^ w46775;
	assign w29951 = w46780 ^ w29827;
	assign w29828 = w29868 ^ w29866;
	assign w29937 = w46780 & w29951;
	assign w49807 = w8951 ^ w8952;
	assign w46777 = w49807 ^ w1017;
	assign w29842 = w46777 ^ w46778;
	assign w29865 = w46779 ^ w46777;
	assign w29944 = w29865 ^ w29828;
	assign w29931 = w29953 & w29944;
	assign w29867 = w46778 ^ w29865;
	assign w29942 = w29872 ^ w29867;
	assign w29943 = w46774 ^ w29867;
	assign w29956 = w46778 ^ w46776;
	assign w29941 = w29866 ^ w29956;
	assign w29932 = w29956 & w29941;
	assign w29934 = w29949 & w29942;
	assign w29940 = w46775 ^ w29867;
	assign w29936 = w29955 & w29940;
	assign w29870 = w29936 ^ w29866;
	assign w44620 = w29931 ^ w29937;
	assign w29881 = w44620 ^ w29866;
	assign w44621 = w29931 ^ w29934;
	assign w29884 = w29932 ^ w44621;
	assign w29844 = w29870 ^ w44621;
	assign w29948 = w46779 ^ w29952;
	assign w29935 = w29952 & w29948;
	assign w29840 = w29935 ^ w29884;
	assign w29922 = w46779 ^ w29840;
	assign w29954 = w46776 ^ w46773;
	assign w29950 = w29954 ^ w29882;
	assign w29933 = w29954 & w29943;
	assign w29841 = w29932 ^ w29933;
	assign w29888 = w29841 ^ w29842;
	assign w29887 = w29888 ^ w29870;
	assign w29929 = w29935 ^ w29887;
	assign w29869 = w29933 ^ w29867;
	assign w29928 = w29844 ^ w29869;
	assign w29946 = w29865 ^ w29954;
	assign w29939 = w29946 & w29950;
	assign w29871 = w29939 ^ w29868;
	assign w29945 = w46780 ^ w29946;
	assign w29938 = w29947 & w29945;
	assign w29889 = w29932 ^ w29938;
	assign w29927 = w29889 ^ w29881;
	assign w29875 = w29871 ^ w29869;
	assign w29843 = w29875 ^ w44620;
	assign w29886 = w46775 ^ w29843;
	assign w29880 = w46773 ^ w29875;
	assign w29930 = w29889 ^ w29880;
	assign w29926 = w29930 & w29929;
	assign w29925 = w29926 ^ w29928;
	assign w29924 = w29927 & w29925;
	assign w29835 = w29924 ^ w29936;
	assign w29832 = w29924 ^ w29880;
	assign w29831 = w29835 ^ w29871;
	assign w29834 = w46773 ^ w29831;
	assign w29830 = w46775 ^ w29831;
	assign w29923 = w29924 ^ w29886;
	assign w29893 = w29923 & w29949;
	assign w29902 = w29923 & w29942;
	assign w29921 = w29926 ^ w29886;
	assign w29920 = w29921 & w29922;
	assign w29839 = w29920 ^ w29884;
	assign w29918 = w29926 ^ w29920;
	assign w29917 = w29928 & w29918;
	assign w29838 = w29920 ^ w29937;
	assign w29833 = w29838 ^ w29934;
	assign w29911 = w29833 ^ w29834;
	assign w29901 = w29911 & w29943;
	assign w29919 = w29920 ^ w29928;
	assign w29905 = w29919 & w46780;
	assign w29896 = w29919 & w29951;
	assign w29915 = w29917 ^ w29925;
	assign w29914 = w29923 & w29915;
	assign w29837 = w29914 ^ w29938;
	assign w29879 = w29914 ^ w29889;
	assign w29910 = w29879 ^ w29832;
	assign w29895 = w29910 & w29955;
	assign w29904 = w29910 & w29940;
	assign w29862 = w29904 ^ w29895;
	assign w29913 = w29879 ^ w29881;
	assign w29903 = w29913 & w29952;
	assign w29846 = w29902 ^ w29903;
	assign w29894 = w29913 & w29948;
	assign w29892 = w29911 & w29954;
	assign w44623 = w29903 ^ w29904;
	assign w44625 = w29917 ^ w29935;
	assign w29909 = w44625 ^ w29887;
	assign w29898 = w29909 & w29950;
	assign w29907 = w29909 & w29946;
	assign w44624 = w29905 ^ w29907;
	assign w29864 = w29902 ^ w29894;
	assign w29876 = w46779 ^ w44625;
	assign w29916 = w29876 ^ w29839;
	assign w29906 = w29916 & w29945;
	assign w29897 = w29916 & w29947;
	assign w29829 = w29876 ^ w29837;
	assign w29836 = w29866 ^ w29829;
	assign w29912 = w29833 ^ w29836;
	assign w29899 = w29912 & w29944;
	assign w29890 = w29912 & w29953;
	assign w29856 = w29901 ^ w29890;
	assign w29908 = w29829 ^ w29830;
	assign w29891 = w29908 & w29956;
	assign w29900 = w29908 & w29941;
	assign w29857 = w29900 ^ w29901;
	assign w29885 = w29900 ^ w44623;
	assign w29851 = w29896 ^ w29885;
	assign w29848 = ~w29851;
	assign w29845 = w29901 ^ w29885;
	assign w29861 = w29900 ^ w29903;
	assign w29852 = ~w29856;
	assign w44622 = w29891 ^ w29892;
	assign w29873 = w29897 ^ w44622;
	assign w29874 = w29898 ^ w29873;
	assign w29878 = w29906 ^ w29874;
	assign w29883 = w29907 ^ w29878;
	assign w29958 = w29883 ^ w29857;
	assign w50099 = w44623 ^ w29883;
	assign w9511 = w50095 ^ w50099;
	assign w9321 = w9298 ^ w9511;
	assign w49993 = w9321 ^ w9322;
	assign w46664 = w49993 ^ w1130;
	assign w9292 = w9516 ^ w9511;
	assign w50010 = w45604 ^ w9292;
	assign w46647 = w50010 ^ w1147;
	assign w9269 = w9268 ^ w50099;
	assign w9557 = w9269 ^ w9270;
	assign w50001 = w9557 ^ w9523;
	assign w46656 = w50001 ^ w1138;
	assign w29847 = w29905 ^ w29878;
	assign w50098 = w29846 ^ w29847;
	assign w9265 = w9268 ^ w50098;
	assign w9558 = w9265 ^ w9266;
	assign w50000 = w9558 ^ w9531;
	assign w9520 = w50094 ^ w50098;
	assign w9293 = w9295 ^ w9520;
	assign w9323 = w9314 ^ w9520;
	assign w49992 = w9323 ^ w9324;
	assign w46657 = w50000 ^ w1137;
	assign w46665 = w49992 ^ w1129;
	assign w29860 = w29864 ^ w44622;
	assign w29863 = w44624 ^ w29860;
	assign w29858 = ~w29861;
	assign w50100 = w29874 ^ w29845;
	assign w9305 = w45896 ^ w50100;
	assign w50004 = w9305 ^ w9306;
	assign w46653 = w50004 ^ w1141;
	assign w15348 = w46656 ^ w46653;
	assign w9488 = w50085 ^ w50100;
	assign w9261 = w9488 ^ w50098;
	assign w9560 = w9261 ^ w9262;
	assign w9257 = ~w9488;
	assign w49985 = w9560 ^ w9511;
	assign w46672 = w49985 ^ w1122;
	assign w9480 = w50096 ^ w50100;
	assign w9318 = w9509 ^ w9480;
	assign w49996 = w50085 ^ w9318;
	assign w9304 = w9546 ^ w9480;
	assign w46661 = w49996 ^ w1133;
	assign w11328 = w46664 ^ w46661;
	assign w50005 = w45599 ^ w9304;
	assign w46652 = w50005 ^ w1142;
	assign w29877 = w29895 ^ w29899;
	assign w29855 = ~w29877;
	assign w29859 = w29855 ^ w29860;
	assign w29959 = w29858 ^ w29859;
	assign w29854 = w29855 ^ w29893;
	assign w29850 = w29854 ^ w44624;
	assign w29849 = w29873 ^ w29850;
	assign w50097 = w29848 ^ w29849;
	assign w9258 = w9257 ^ w50097;
	assign w9530 = w50093 ^ w50097;
	assign w9296 = w9298 ^ w9530;
	assign w9561 = w9258 ^ w9259;
	assign w49984 = w9561 ^ w9520;
	assign w46673 = w49984 ^ w1121;
	assign w29853 = w29892 ^ w29850;
	assign w29957 = w29852 ^ w29853;
	assign w9312 = w9314 ^ w50097;
	assign w49999 = w9312 ^ w9313;
	assign w46658 = w49999 ^ w1136;
	assign w15236 = w46657 ^ w46658;
	assign w15347 = w46653 ^ w46658;
	assign w15350 = w46658 ^ w46656;
	assign w29960 = w29862 ^ w29863;
	assign w9343 = ~w9530;
	assign w9325 = w9545 ^ w9530;
	assign w49991 = w50082 ^ w9325;
	assign w46666 = w49991 ^ w1128;
	assign w11327 = w46661 ^ w46666;
	assign w11330 = w46666 ^ w46664;
	assign w45682 = ~w29957;
	assign w9310 = w9516 ^ w45682;
	assign w9505 = w45604 ^ w45682;
	assign w9320 = w9523 ^ w9505;
	assign w9291 = w9509 ^ w9505;
	assign w50011 = w45605 ^ w9291;
	assign w46646 = w50011 ^ w1148;
	assign w23708 = w46652 ^ w46646;
	assign w23788 = w46647 ^ w23708;
	assign w9340 = w9505 ^ w50099;
	assign w9338 = ~w9340;
	assign w49986 = w9338 ^ w9339;
	assign w46671 = w49986 ^ w1123;
	assign w49994 = w45600 ^ w9320;
	assign w46663 = w49994 ^ w1131;
	assign w11240 = w46663 ^ w46661;
	assign w11315 = w11240 ^ w11330;
	assign w50002 = w9310 ^ w9311;
	assign w46655 = w50002 ^ w1139;
	assign w15260 = w46655 ^ w46653;
	assign w15335 = w15260 ^ w15350;
	assign w15326 = w15350 & w15335;
	assign w11306 = w11330 & w11315;
	assign w45683 = ~w29958;
	assign w9330 = w9480 ^ w45683;
	assign w49988 = w9330 ^ w9331;
	assign w46669 = w49988 ^ w1125;
	assign w26604 = w46672 ^ w46669;
	assign w26516 = w46671 ^ w46669;
	assign w9494 = w45605 ^ w45683;
	assign w9333 = w9494 ^ w45682;
	assign w9319 = w9516 ^ w9494;
	assign w49995 = w45601 ^ w9319;
	assign w9290 = w9494 ^ w9483;
	assign w50012 = w50096 ^ w9290;
	assign w46645 = w50012 ^ w1149;
	assign w46662 = w49995 ^ w1132;
	assign w11242 = w46664 ^ w46662;
	assign w11202 = w11242 ^ w11240;
	assign w11201 = w11242 ^ w46663;
	assign w23702 = w46647 ^ w46645;
	assign w23785 = w23702 ^ w23708;
	assign w9332 = w9333 ^ w9334;
	assign w49987 = ~w9332;
	assign w46670 = w49987 ^ w1124;
	assign w26518 = w46672 ^ w46670;
	assign w26477 = w26518 ^ w46671;
	assign w26478 = w26518 ^ w26516;
	assign w45684 = ~w29959;
	assign w9341 = w9343 ^ w45684;
	assign w49983 = w9341 ^ w9342;
	assign w9534 = w45598 ^ w45684;
	assign w9299 = w9538 ^ w9534;
	assign w50007 = w50093 ^ w9299;
	assign w9327 = w9546 ^ w9534;
	assign w9326 = w9327 ^ w9328;
	assign w46674 = w49983 ^ w1120;
	assign w26492 = w46673 ^ w46674;
	assign w26606 = w46674 ^ w46672;
	assign w26591 = w26516 ^ w26606;
	assign w26603 = w46669 ^ w46674;
	assign w46650 = w50007 ^ w1144;
	assign w23789 = w46645 ^ w46650;
	assign w26582 = w26606 & w26591;
	assign w49990 = ~w9326;
	assign w46667 = w49990 ^ w1127;
	assign w11239 = w46667 ^ w46665;
	assign w11318 = w11239 ^ w11202;
	assign w11305 = w11327 & w11318;
	assign w11329 = w46661 ^ w46667;
	assign w11256 = w46667 ^ w46666;
	assign w11324 = w11328 ^ w11256;
	assign w11241 = w46666 ^ w11239;
	assign w11317 = w46662 ^ w11241;
	assign w11307 = w11328 & w11317;
	assign w11243 = w11307 ^ w11241;
	assign w11215 = w11306 ^ w11307;
	assign w11314 = w46663 ^ w11241;
	assign w11310 = w11329 & w11314;
	assign w11244 = w11310 ^ w11240;
	assign w11320 = w11239 ^ w11328;
	assign w11313 = w11320 & w11324;
	assign w9263 = w9487 ^ w45684;
	assign w9559 = w9263 ^ w9264;
	assign w49998 = w9559 ^ w9545;
	assign w46659 = w49998 ^ w1135;
	assign w15349 = w46653 ^ w46659;
	assign w15259 = w46659 ^ w46657;
	assign w15340 = w15259 ^ w15348;
	assign w15261 = w46658 ^ w15259;
	assign w15334 = w46655 ^ w15261;
	assign w15330 = w15349 & w15334;
	assign w15264 = w15330 ^ w15260;
	assign w15276 = w46659 ^ w46658;
	assign w15344 = w15348 ^ w15276;
	assign w15333 = w15340 & w15344;
	assign w11245 = w11313 ^ w11242;
	assign w11249 = w11245 ^ w11243;
	assign w11254 = w46661 ^ w11249;
	assign w45685 = ~w29960;
	assign w9255 = w9257 ^ w45685;
	assign w49997 = w45685 ^ w9315;
	assign w9542 = w45599 ^ w45685;
	assign w9303 = w9545 ^ w9542;
	assign w9329 = w9542 ^ w9483;
	assign w49989 = w45595 ^ w9329;
	assign w46668 = w49989 ^ w1126;
	assign w11325 = w46668 ^ w11201;
	assign w11311 = w46668 & w11325;
	assign w11246 = w46668 ^ w46662;
	assign w11316 = w11246 ^ w11241;
	assign w11323 = w11240 ^ w11246;
	assign w11321 = w11256 ^ w11323;
	assign w11326 = w46663 ^ w11246;
	assign w11322 = w46667 ^ w11326;
	assign w11319 = w46668 ^ w11320;
	assign w11312 = w11321 & w11319;
	assign w11309 = w11326 & w11322;
	assign w46660 = w49997 ^ w1134;
	assign w15339 = w46660 ^ w15340;
	assign w9562 = w9255 ^ w9256;
	assign w49982 = w9562 ^ w9534;
	assign w46675 = w49982 ^ w1119;
	assign w26532 = w46675 ^ w46674;
	assign w26605 = w46669 ^ w46675;
	assign w26600 = w26604 ^ w26532;
	assign w26515 = w46675 ^ w46673;
	assign w26596 = w26515 ^ w26604;
	assign w26589 = w26596 & w26600;
	assign w26517 = w46674 ^ w26515;
	assign w26593 = w46670 ^ w26517;
	assign w26583 = w26604 & w26593;
	assign w26519 = w26583 ^ w26517;
	assign w43845 = w11305 ^ w11311;
	assign w11217 = w11249 ^ w43845;
	assign w11255 = w43845 ^ w11240;
	assign w26521 = w26589 ^ w26518;
	assign w26525 = w26521 ^ w26519;
	assign w26530 = w46669 ^ w26525;
	assign w11308 = w11323 & w11316;
	assign w43842 = w11305 ^ w11308;
	assign w26491 = w26582 ^ w26583;
	assign w26538 = w26491 ^ w26492;
	assign w11258 = w11306 ^ w43842;
	assign w26594 = w26515 ^ w26478;
	assign w26581 = w26603 & w26594;
	assign w9301 = ~w9303;
	assign w9344 = w9542 ^ w9488;
	assign w49981 = w45234 ^ w9344;
	assign w46676 = w49981 ^ w1118;
	assign w26522 = w46676 ^ w46670;
	assign w26599 = w26516 ^ w26522;
	assign w26595 = w46676 ^ w26596;
	assign w26592 = w26522 ^ w26517;
	assign w26601 = w46676 ^ w26477;
	assign w26602 = w46671 ^ w26522;
	assign w26598 = w46675 ^ w26602;
	assign w26597 = w26532 ^ w26599;
	assign w26588 = w26597 & w26595;
	assign w26585 = w26602 & w26598;
	assign w26587 = w46676 & w26601;
	assign w26539 = w26582 ^ w26588;
	assign w26580 = w26539 ^ w26530;
	assign w44482 = w26581 ^ w26587;
	assign w26493 = w26525 ^ w44482;
	assign w26536 = w46671 ^ w26493;
	assign w26531 = w44482 ^ w26516;
	assign w26577 = w26539 ^ w26531;
	assign w26584 = w26599 & w26592;
	assign w44479 = w26581 ^ w26584;
	assign w26534 = w26582 ^ w44479;
	assign w26490 = w26585 ^ w26534;
	assign w11263 = w11306 ^ w11312;
	assign w11304 = w11263 ^ w11254;
	assign w11301 = w11263 ^ w11255;
	assign w26590 = w46671 ^ w26517;
	assign w26586 = w26605 & w26590;
	assign w26520 = w26586 ^ w26516;
	assign w26537 = w26538 ^ w26520;
	assign w26579 = w26585 ^ w26537;
	assign w26576 = w26580 & w26579;
	assign w26571 = w26576 ^ w26536;
	assign w26494 = w26520 ^ w44479;
	assign w26578 = w26494 ^ w26519;
	assign w26575 = w26576 ^ w26578;
	assign w26574 = w26577 & w26575;
	assign w26573 = w26574 ^ w26536;
	assign w26543 = w26573 & w26599;
	assign w26485 = w26574 ^ w26586;
	assign w26481 = w26485 ^ w26521;
	assign w26484 = w46669 ^ w26481;
	assign w26482 = w26574 ^ w26530;
	assign w26552 = w26573 & w26592;
	assign w26480 = w46671 ^ w26481;
	assign w11218 = w11244 ^ w43842;
	assign w11302 = w11218 ^ w11243;
	assign w11260 = w46663 ^ w11217;
	assign w11216 = w46665 ^ w46666;
	assign w11262 = w11215 ^ w11216;
	assign w11261 = w11262 ^ w11244;
	assign w11303 = w11309 ^ w11261;
	assign w11300 = w11304 & w11303;
	assign w11299 = w11300 ^ w11302;
	assign w11298 = w11301 & w11299;
	assign w11209 = w11298 ^ w11310;
	assign w11297 = w11298 ^ w11260;
	assign w11276 = w11297 & w11316;
	assign w11206 = w11298 ^ w11254;
	assign w11205 = w11209 ^ w11245;
	assign w11208 = w46661 ^ w11205;
	assign w11204 = w46663 ^ w11205;
	assign w11267 = w11297 & w11323;
	assign w11295 = w11300 ^ w11260;
	assign w11214 = w11309 ^ w11258;
	assign w11296 = w46667 ^ w11214;
	assign w11294 = w11295 & w11296;
	assign w11293 = w11294 ^ w11302;
	assign w11270 = w11293 & w11325;
	assign w11279 = w11293 & w46668;
	assign w11213 = w11294 ^ w11258;
	assign w11292 = w11300 ^ w11294;
	assign w11291 = w11302 & w11292;
	assign w11289 = w11291 ^ w11299;
	assign w43844 = w11291 ^ w11309;
	assign w11288 = w11297 & w11289;
	assign w11253 = w11288 ^ w11263;
	assign w11284 = w11253 ^ w11206;
	assign w11269 = w11284 & w11329;
	assign w11278 = w11284 & w11314;
	assign w11236 = w11278 ^ w11269;
	assign w11211 = w11288 ^ w11312;
	assign w11283 = w43844 ^ w11261;
	assign w11281 = w11283 & w11320;
	assign w43847 = w11279 ^ w11281;
	assign w11272 = w11283 & w11324;
	assign w11250 = w46667 ^ w43844;
	assign w11203 = w11250 ^ w11211;
	assign w11282 = w11203 ^ w11204;
	assign w11265 = w11282 & w11330;
	assign w11274 = w11282 & w11315;
	assign w11210 = w11240 ^ w11203;
	assign w11290 = w11250 ^ w11213;
	assign w11271 = w11290 & w11321;
	assign w11280 = w11290 & w11319;
	assign w11287 = w11253 ^ w11255;
	assign w11277 = w11287 & w11326;
	assign w11220 = w11276 ^ w11277;
	assign w11235 = w11274 ^ w11277;
	assign w11268 = w11287 & w11322;
	assign w11238 = w11276 ^ w11268;
	assign w43846 = w11277 ^ w11278;
	assign w11259 = w11274 ^ w43846;
	assign w11232 = ~w11235;
	assign w11225 = w11270 ^ w11259;
	assign w11222 = ~w11225;
	assign w11212 = w11294 ^ w11311;
	assign w11207 = w11212 ^ w11308;
	assign w11286 = w11207 ^ w11210;
	assign w11273 = w11286 & w11318;
	assign w11251 = w11269 ^ w11273;
	assign w11285 = w11207 ^ w11208;
	assign w11266 = w11285 & w11328;
	assign w11229 = ~w11251;
	assign w11264 = w11286 & w11327;
	assign w11275 = w11285 & w11317;
	assign w11230 = w11275 ^ w11264;
	assign w11219 = w11275 ^ w11259;
	assign w11226 = ~w11230;
	assign w11231 = w11274 ^ w11275;
	assign w11228 = w11229 ^ w11267;
	assign w11224 = w11228 ^ w43847;
	assign w11227 = w11266 ^ w11224;
	assign w11331 = w11226 ^ w11227;
	assign w50253 = ~w11331;
	assign w43476 = w45324 ^ w50253;
	assign w43351 = w45588 ^ w11331;
	assign w43843 = w11265 ^ w11266;
	assign w11234 = w11238 ^ w43843;
	assign w11237 = w43847 ^ w11234;
	assign w11334 = w11236 ^ w11237;
	assign w11233 = w11229 ^ w11234;
	assign w11333 = w11232 ^ w11233;
	assign w45227 = ~w11333;
	assign w43465 = w45227 ^ w50256;
	assign w45228 = ~w11334;
	assign w43464 = w45228 ^ w45582;
	assign w11247 = w11271 ^ w43843;
	assign w11223 = w11247 ^ w11224;
	assign w50250 = w11222 ^ w11223;
	assign w43463 = w50250 ^ w50257;
	assign w43346 = ~w43463;
	assign w43344 = w43346 ^ w50246;
	assign w43215 = w50246 ^ w50250;
	assign w11248 = w11272 ^ w11247;
	assign w11252 = w11280 ^ w11248;
	assign w11221 = w11279 ^ w11252;
	assign w50255 = w11248 ^ w11219;
	assign w11257 = w11281 ^ w11252;
	assign w50252 = w43846 ^ w11257;
	assign w43424 = w50249 ^ w50255;
	assign w43425 = w50255 ^ w50260;
	assign w43479 = w50248 ^ w50252;
	assign w43359 = ~w43425;
	assign w43363 = w43359 ^ w45227;
	assign w43353 = w50259 ^ w50252;
	assign w43214 = w43424 ^ w50247;
	assign w43493 = w43214 ^ w43215;
	assign w11332 = w11257 ^ w11231;
	assign w50254 = ~w11332;
	assign w43474 = w45325 ^ w50254;
	assign w43349 = w45589 ^ w11332;
	assign w50251 = w11220 ^ w11221;
	assign w43488 = w50247 ^ w50251;
	assign w43370 = ~w43488;
	assign w43357 = w43488 ^ w43346;
	assign w43211 = w50258 ^ w50251;
	assign w9309 = w9509 ^ w45683;
	assign w9307 = ~w9309;
	assign w50003 = w9307 ^ w9308;
	assign w46654 = w50003 ^ w1140;
	assign w15266 = w46660 ^ w46654;
	assign w15336 = w15266 ^ w15261;
	assign w15346 = w46655 ^ w15266;
	assign w15337 = w46654 ^ w15261;
	assign w15327 = w15348 & w15337;
	assign w15235 = w15326 ^ w15327;
	assign w15263 = w15327 ^ w15261;
	assign w15282 = w15235 ^ w15236;
	assign w15281 = w15282 ^ w15264;
	assign w15343 = w15260 ^ w15266;
	assign w15328 = w15343 & w15336;
	assign w15262 = w46656 ^ w46654;
	assign w15222 = w15262 ^ w15260;
	assign w15338 = w15259 ^ w15222;
	assign w15221 = w15262 ^ w46655;
	assign w15325 = w15347 & w15338;
	assign w15345 = w46660 ^ w15221;
	assign w15331 = w46660 & w15345;
	assign w15265 = w15333 ^ w15262;
	assign w15269 = w15265 ^ w15263;
	assign w15274 = w46653 ^ w15269;
	assign w15341 = w15276 ^ w15343;
	assign w15332 = w15341 & w15339;
	assign w15342 = w46659 ^ w15346;
	assign w15329 = w15346 & w15342;
	assign w15323 = w15329 ^ w15281;
	assign w44008 = w15325 ^ w15331;
	assign w15237 = w15269 ^ w44008;
	assign w15280 = w46655 ^ w15237;
	assign w15275 = w44008 ^ w15260;
	assign w44009 = w15325 ^ w15328;
	assign w15278 = w15326 ^ w44009;
	assign w15234 = w15329 ^ w15278;
	assign w15316 = w46659 ^ w15234;
	assign w15238 = w15264 ^ w44009;
	assign w15322 = w15238 ^ w15263;
	assign w15283 = w15326 ^ w15332;
	assign w15324 = w15283 ^ w15274;
	assign w15320 = w15324 & w15323;
	assign w15315 = w15320 ^ w15280;
	assign w15314 = w15315 & w15316;
	assign w15313 = w15314 ^ w15322;
	assign w15312 = w15320 ^ w15314;
	assign w15311 = w15322 & w15312;
	assign w15233 = w15314 ^ w15278;
	assign w15232 = w15314 ^ w15331;
	assign w15227 = w15232 ^ w15328;
	assign w15319 = w15320 ^ w15322;
	assign w15309 = w15311 ^ w15319;
	assign w15299 = w15313 & w46660;
	assign w15290 = w15313 & w15345;
	assign w15321 = w15283 ^ w15275;
	assign w15318 = w15321 & w15319;
	assign w15226 = w15318 ^ w15274;
	assign w15317 = w15318 ^ w15280;
	assign w15296 = w15317 & w15336;
	assign w15287 = w15317 & w15343;
	assign w15308 = w15317 & w15309;
	assign w15231 = w15308 ^ w15332;
	assign w15229 = w15318 ^ w15330;
	assign w15225 = w15229 ^ w15265;
	assign w15228 = w46653 ^ w15225;
	assign w15305 = w15227 ^ w15228;
	assign w15295 = w15305 & w15337;
	assign w15286 = w15305 & w15348;
	assign w15224 = w46655 ^ w15225;
	assign w15273 = w15308 ^ w15283;
	assign w15307 = w15273 ^ w15275;
	assign w15304 = w15273 ^ w15226;
	assign w15298 = w15304 & w15334;
	assign w15288 = w15307 & w15342;
	assign w15297 = w15307 & w15346;
	assign w15240 = w15296 ^ w15297;
	assign w15289 = w15304 & w15349;
	assign w15256 = w15298 ^ w15289;
	assign w44011 = w15297 ^ w15298;
	assign w15258 = w15296 ^ w15288;
	assign w44013 = w15311 ^ w15329;
	assign w15270 = w46659 ^ w44013;
	assign w15223 = w15270 ^ w15231;
	assign w15302 = w15223 ^ w15224;
	assign w15294 = w15302 & w15335;
	assign w15251 = w15294 ^ w15295;
	assign w15285 = w15302 & w15350;
	assign w15230 = w15260 ^ w15223;
	assign w15306 = w15227 ^ w15230;
	assign w15293 = w15306 & w15338;
	assign w15284 = w15306 & w15347;
	assign w15310 = w15270 ^ w15233;
	assign w15300 = w15310 & w15339;
	assign w15291 = w15310 & w15341;
	assign w15271 = w15289 ^ w15293;
	assign w15249 = ~w15271;
	assign w15248 = w15249 ^ w15287;
	assign w15279 = w15294 ^ w44011;
	assign w15239 = w15295 ^ w15279;
	assign w15245 = w15290 ^ w15279;
	assign w15242 = ~w15245;
	assign w44010 = w15285 ^ w15286;
	assign w15267 = w15291 ^ w44010;
	assign w15254 = w15258 ^ w44010;
	assign w15253 = w15249 ^ w15254;
	assign w15255 = w15294 ^ w15297;
	assign w15252 = ~w15255;
	assign w15353 = w15252 ^ w15253;
	assign w15250 = w15295 ^ w15284;
	assign w15246 = ~w15250;
	assign w15303 = w44013 ^ w15281;
	assign w15292 = w15303 & w15344;
	assign w15301 = w15303 & w15340;
	assign w44012 = w15299 ^ w15301;
	assign w15244 = w15248 ^ w44012;
	assign w15247 = w15286 ^ w15244;
	assign w15243 = w15267 ^ w15244;
	assign w50311 = w15242 ^ w15243;
	assign w15351 = w15246 ^ w15247;
	assign w15268 = w15292 ^ w15267;
	assign w50314 = w15268 ^ w15239;
	assign w15272 = w15300 ^ w15268;
	assign w15241 = w15299 ^ w15272;
	assign w50312 = w15240 ^ w15241;
	assign w15277 = w15301 ^ w15272;
	assign w50313 = w44011 ^ w15277;
	assign w15352 = w15277 ^ w15251;
	assign w43225 = w50313 ^ w50312;
	assign w15257 = w44012 ^ w15254;
	assign w15354 = w15256 ^ w15257;
	assign w45310 = ~w15353;
	assign w45311 = ~w15354;
	assign w45316 = ~w15351;
	assign w45317 = ~w15352;
	assign w43373 = w45317 ^ w45316;
	assign w26572 = w46675 ^ w26490;
	assign w26570 = w26571 & w26572;
	assign w26569 = w26570 ^ w26578;
	assign w26546 = w26569 & w26601;
	assign w26568 = w26576 ^ w26570;
	assign w26488 = w26570 ^ w26587;
	assign w26483 = w26488 ^ w26584;
	assign w26561 = w26483 ^ w26484;
	assign w26551 = w26561 & w26593;
	assign w26542 = w26561 & w26604;
	assign w26567 = w26578 & w26568;
	assign w26565 = w26567 ^ w26575;
	assign w26564 = w26573 & w26565;
	assign w26487 = w26564 ^ w26588;
	assign w44481 = w26567 ^ w26585;
	assign w26559 = w44481 ^ w26537;
	assign w26526 = w46675 ^ w44481;
	assign w26479 = w26526 ^ w26487;
	assign w26558 = w26479 ^ w26480;
	assign w26550 = w26558 & w26591;
	assign w26486 = w26516 ^ w26479;
	assign w26562 = w26483 ^ w26486;
	assign w26541 = w26558 & w26606;
	assign w26540 = w26562 & w26603;
	assign w26506 = w26551 ^ w26540;
	assign w26502 = ~w26506;
	assign w44480 = w26541 ^ w26542;
	assign w26529 = w26564 ^ w26539;
	assign w26563 = w26529 ^ w26531;
	assign w26544 = w26563 & w26598;
	assign w26553 = w26563 & w26602;
	assign w26496 = w26552 ^ w26553;
	assign w26511 = w26550 ^ w26553;
	assign w26508 = ~w26511;
	assign w26514 = w26552 ^ w26544;
	assign w26510 = w26514 ^ w44480;
	assign w26560 = w26529 ^ w26482;
	assign w26545 = w26560 & w26605;
	assign w26554 = w26560 & w26590;
	assign w26512 = w26554 ^ w26545;
	assign w44483 = w26553 ^ w26554;
	assign w26535 = w26550 ^ w44483;
	assign w26501 = w26546 ^ w26535;
	assign w26498 = ~w26501;
	assign w26495 = w26551 ^ w26535;
	assign w26557 = w26559 & w26596;
	assign w26549 = w26562 & w26594;
	assign w26527 = w26545 ^ w26549;
	assign w26505 = ~w26527;
	assign w26509 = w26505 ^ w26510;
	assign w26504 = w26505 ^ w26543;
	assign w26609 = w26508 ^ w26509;
	assign w45586 = ~w26609;
	assign w26555 = w26569 & w46676;
	assign w44484 = w26555 ^ w26557;
	assign w26513 = w44484 ^ w26510;
	assign w26610 = w26512 ^ w26513;
	assign w26500 = w26504 ^ w44484;
	assign w26503 = w26542 ^ w26500;
	assign w26607 = w26502 ^ w26503;
	assign w45587 = ~w26610;
	assign w45592 = ~w26607;
	assign w43331 = w45681 ^ w45592;
	assign w26507 = w26550 ^ w26551;
	assign w26548 = w26559 & w26600;
	assign w26489 = w26570 ^ w26534;
	assign w26566 = w26526 ^ w26489;
	assign w26556 = w26566 & w26595;
	assign w26547 = w26566 & w26597;
	assign w26523 = w26547 ^ w44480;
	assign w26499 = w26523 ^ w26500;
	assign w26524 = w26548 ^ w26523;
	assign w50269 = w26524 ^ w26495;
	assign w26528 = w26556 ^ w26524;
	assign w26533 = w26557 ^ w26528;
	assign w50268 = w44483 ^ w26533;
	assign w26608 = w26533 ^ w26507;
	assign w43430 = w50269 ^ w50282;
	assign w43181 = w43430 ^ w50280;
	assign w43177 = ~w43430;
	assign w43178 = w43177 ^ w50279;
	assign w43175 = w43177 ^ w45676;
	assign w50266 = w26498 ^ w26499;
	assign w45593 = ~w26608;
	assign w43439 = w45593 ^ w45674;
	assign w43312 = w50269 ^ w45593;
	assign w26497 = w26555 ^ w26528;
	assign w50267 = w26496 ^ w26497;
	assign w45944 = ~w9478;
	assign w9441 = w45944 ^ w45332;
	assign w9469 = w45944 ^ w45514;
	assign w50020 = w9469 ^ w9470;
	assign w50038 = w9440 ^ w9441;
	assign w9438 = w45944 ^ w50102;
	assign w9436 = w9437 ^ w9438;
	assign w50040 = ~w9436;
	assign w46617 = w50040 ^ w1113;
	assign w29440 = w46617 ^ w46618;
	assign w46619 = w50038 ^ w1111;
	assign w29480 = w46619 ^ w46618;
	assign w29548 = w29552 ^ w29480;
	assign w29553 = w46613 ^ w46619;
	assign w29545 = w29480 ^ w29547;
	assign w46637 = w50020 ^ w1093;
	assign w15126 = w46639 ^ w46637;
	assign w15201 = w15126 ^ w15216;
	assign w15209 = w15126 ^ w15132;
	assign w15214 = w46640 ^ w46637;
	assign w15206 = w15125 ^ w15214;
	assign w15205 = w46644 ^ w15206;
	assign w15193 = w15214 & w15203;
	assign w15129 = w15193 ^ w15127;
	assign w15210 = w15214 ^ w15142;
	assign w15207 = w15142 ^ w15209;
	assign w15198 = w15207 & w15205;
	assign w29546 = w46619 ^ w29550;
	assign w29463 = w46619 ^ w46617;
	assign w29544 = w29463 ^ w29552;
	assign w29543 = w46620 ^ w29544;
	assign w29465 = w46618 ^ w29463;
	assign w29538 = w46615 ^ w29465;
	assign w29541 = w46614 ^ w29465;
	assign w29531 = w29552 & w29541;
	assign w29439 = w29530 ^ w29531;
	assign w29486 = w29439 ^ w29440;
	assign w29467 = w29531 ^ w29465;
	assign w29540 = w29470 ^ w29465;
	assign w29532 = w29547 & w29540;
	assign w29537 = w29544 & w29548;
	assign w29469 = w29537 ^ w29466;
	assign w29473 = w29469 ^ w29467;
	assign w29478 = w46613 ^ w29473;
	assign w29536 = w29545 & w29543;
	assign w29487 = w29530 ^ w29536;
	assign w29528 = w29487 ^ w29478;
	assign w29542 = w29463 ^ w29426;
	assign w29529 = w29551 & w29542;
	assign w44603 = w29529 ^ w29535;
	assign w29441 = w29473 ^ w44603;
	assign w29479 = w44603 ^ w29464;
	assign w29525 = w29487 ^ w29479;
	assign w44604 = w29529 ^ w29532;
	assign w29482 = w29530 ^ w44604;
	assign w29484 = w46615 ^ w29441;
	assign w29533 = w29550 & w29546;
	assign w29438 = w29533 ^ w29482;
	assign w29520 = w46619 ^ w29438;
	assign w15088 = w15128 ^ w15126;
	assign w15204 = w15125 ^ w15088;
	assign w15215 = w46637 ^ w46643;
	assign w15213 = w46637 ^ w46642;
	assign w15199 = w15206 & w15210;
	assign w15131 = w15199 ^ w15128;
	assign w15135 = w15131 ^ w15129;
	assign w15140 = w46637 ^ w15135;
	assign w15196 = w15215 & w15200;
	assign w15130 = w15196 ^ w15126;
	assign w15194 = w15209 & w15202;
	assign w15192 = w15216 & w15201;
	assign w15149 = w15192 ^ w15198;
	assign w15190 = w15149 ^ w15140;
	assign w15191 = w15213 & w15204;
	assign w44003 = w15191 ^ w15197;
	assign w15141 = w44003 ^ w15126;
	assign w15187 = w15149 ^ w15141;
	assign w15103 = w15135 ^ w44003;
	assign w44004 = w15191 ^ w15194;
	assign w15144 = w15192 ^ w44004;
	assign w15100 = w15195 ^ w15144;
	assign w15182 = w46643 ^ w15100;
	assign w15104 = w15130 ^ w44004;
	assign w15188 = w15104 ^ w15129;
	assign w15146 = w46639 ^ w15103;
	assign w15101 = w15192 ^ w15193;
	assign w15148 = w15101 ^ w15102;
	assign w15147 = w15148 ^ w15130;
	assign w15189 = w15195 ^ w15147;
	assign w15186 = w15190 & w15189;
	assign w15185 = w15186 ^ w15188;
	assign w15181 = w15186 ^ w15146;
	assign w15180 = w15181 & w15182;
	assign w15098 = w15180 ^ w15197;
	assign w15178 = w15186 ^ w15180;
	assign w15099 = w15180 ^ w15144;
	assign w15179 = w15180 ^ w15188;
	assign w15156 = w15179 & w15211;
	assign w15165 = w15179 & w46644;
	assign w15093 = w15098 ^ w15194;
	assign w15184 = w15187 & w15185;
	assign w15183 = w15184 ^ w15146;
	assign w15162 = w15183 & w15202;
	assign w15092 = w15184 ^ w15140;
	assign w15153 = w15183 & w15209;
	assign w15095 = w15184 ^ w15196;
	assign w15091 = w15095 ^ w15131;
	assign w15094 = w46637 ^ w15091;
	assign w15171 = w15093 ^ w15094;
	assign w15152 = w15171 & w15214;
	assign w15161 = w15171 & w15203;
	assign w15090 = w46639 ^ w15091;
	assign w15177 = w15188 & w15178;
	assign w15175 = w15177 ^ w15185;
	assign w15174 = w15183 & w15175;
	assign w15097 = w15174 ^ w15198;
	assign w44007 = w15177 ^ w15195;
	assign w15136 = w46643 ^ w44007;
	assign w15176 = w15136 ^ w15099;
	assign w15089 = w15136 ^ w15097;
	assign w15096 = w15126 ^ w15089;
	assign w15172 = w15093 ^ w15096;
	assign w15159 = w15172 & w15204;
	assign w15150 = w15172 & w15213;
	assign w15116 = w15161 ^ w15150;
	assign w15166 = w15176 & w15205;
	assign w15112 = ~w15116;
	assign w15157 = w15176 & w15207;
	assign w15169 = w44007 ^ w15147;
	assign w15158 = w15169 & w15210;
	assign w15167 = w15169 & w15206;
	assign w44006 = w15165 ^ w15167;
	assign w15139 = w15174 ^ w15149;
	assign w15173 = w15139 ^ w15141;
	assign w15154 = w15173 & w15208;
	assign w15124 = w15162 ^ w15154;
	assign w15163 = w15173 & w15212;
	assign w15106 = w15162 ^ w15163;
	assign w15170 = w15139 ^ w15092;
	assign w15155 = w15170 & w15215;
	assign w15137 = w15155 ^ w15159;
	assign w15115 = ~w15137;
	assign w15114 = w15115 ^ w15153;
	assign w15110 = w15114 ^ w44006;
	assign w15113 = w15152 ^ w15110;
	assign w15217 = w15112 ^ w15113;
	assign w15164 = w15170 & w15200;
	assign w15122 = w15164 ^ w15155;
	assign w44005 = w15163 ^ w15164;
	assign w45312 = ~w15217;
	assign w15168 = w15089 ^ w15090;
	assign w15160 = w15168 & w15201;
	assign w15151 = w15168 & w15216;
	assign w15117 = w15160 ^ w15161;
	assign w15145 = w15160 ^ w44005;
	assign w15111 = w15156 ^ w15145;
	assign w15105 = w15161 ^ w15145;
	assign w15121 = w15160 ^ w15163;
	assign w15118 = ~w15121;
	assign w43540 = w15151 ^ w15152;
	assign w15133 = w15157 ^ w43540;
	assign w15109 = w15133 ^ w15110;
	assign w15108 = ~w15111;
	assign w15134 = w15158 ^ w15133;
	assign w15138 = w15166 ^ w15134;
	assign w15107 = w15165 ^ w15138;
	assign w15143 = w15167 ^ w15138;
	assign w15218 = w15143 ^ w15117;
	assign w50286 = w15134 ^ w15105;
	assign w50284 = w15106 ^ w15107;
	assign w15120 = w15124 ^ w43540;
	assign w15119 = w15115 ^ w15120;
	assign w15219 = w15118 ^ w15119;
	assign w15123 = w44006 ^ w15120;
	assign w15220 = w15122 ^ w15123;
	assign w50285 = w44005 ^ w15143;
	assign w45306 = ~w15219;
	assign w45307 = ~w15220;
	assign w45313 = ~w15218;
	assign w50283 = w15108 ^ w15109;
	assign w29534 = w29553 & w29538;
	assign w29468 = w29534 ^ w29464;
	assign w29485 = w29486 ^ w29468;
	assign w29527 = w29533 ^ w29485;
	assign w29524 = w29528 & w29527;
	assign w29519 = w29524 ^ w29484;
	assign w29518 = w29519 & w29520;
	assign w29436 = w29518 ^ w29535;
	assign w29516 = w29524 ^ w29518;
	assign w29431 = w29436 ^ w29532;
	assign w29437 = w29518 ^ w29482;
	assign w29442 = w29468 ^ w44604;
	assign w29526 = w29442 ^ w29467;
	assign w29515 = w29526 & w29516;
	assign w29523 = w29524 ^ w29526;
	assign w29513 = w29515 ^ w29523;
	assign w29522 = w29525 & w29523;
	assign w29433 = w29522 ^ w29534;
	assign w29521 = w29522 ^ w29484;
	assign w29500 = w29521 & w29540;
	assign w29512 = w29521 & w29513;
	assign w29435 = w29512 ^ w29536;
	assign w29517 = w29518 ^ w29526;
	assign w29494 = w29517 & w29549;
	assign w29429 = w29433 ^ w29469;
	assign w29432 = w46613 ^ w29429;
	assign w29428 = w46615 ^ w29429;
	assign w29503 = w29517 & w46620;
	assign w29477 = w29512 ^ w29487;
	assign w29511 = w29477 ^ w29479;
	assign w29501 = w29511 & w29550;
	assign w29509 = w29431 ^ w29432;
	assign w29490 = w29509 & w29552;
	assign w29499 = w29509 & w29541;
	assign w44608 = w29515 ^ w29533;
	assign w29507 = w44608 ^ w29485;
	assign w29496 = w29507 & w29548;
	assign w29505 = w29507 & w29544;
	assign w44607 = w29503 ^ w29505;
	assign w29474 = w46619 ^ w44608;
	assign w29427 = w29474 ^ w29435;
	assign w29514 = w29474 ^ w29437;
	assign w29504 = w29514 & w29543;
	assign w29495 = w29514 & w29545;
	assign w29434 = w29464 ^ w29427;
	assign w29510 = w29431 ^ w29434;
	assign w29488 = w29510 & w29551;
	assign w29454 = w29499 ^ w29488;
	assign w29497 = w29510 & w29542;
	assign w29430 = w29522 ^ w29478;
	assign w29508 = w29477 ^ w29430;
	assign w29502 = w29508 & w29538;
	assign w29493 = w29508 & w29553;
	assign w29460 = w29502 ^ w29493;
	assign w29475 = w29493 ^ w29497;
	assign w29453 = ~w29475;
	assign w44606 = w29501 ^ w29502;
	assign w29506 = w29427 ^ w29428;
	assign w29498 = w29506 & w29539;
	assign w29483 = w29498 ^ w44606;
	assign w29449 = w29494 ^ w29483;
	assign w29443 = w29499 ^ w29483;
	assign w29489 = w29506 & w29554;
	assign w29459 = w29498 ^ w29501;
	assign w29456 = ~w29459;
	assign w44605 = w29489 ^ w29490;
	assign w29471 = w29495 ^ w44605;
	assign w29472 = w29496 ^ w29471;
	assign w50318 = w29472 ^ w29443;
	assign w43417 = w50314 ^ w50318;
	assign w29476 = w29504 ^ w29472;
	assign w29481 = w29505 ^ w29476;
	assign w50317 = w44606 ^ w29481;
	assign w43434 = w50313 ^ w50317;
	assign w29455 = w29498 ^ w29499;
	assign w29492 = w29511 & w29546;
	assign w29462 = w29500 ^ w29492;
	assign w29458 = w29462 ^ w44605;
	assign w29461 = w44607 ^ w29458;
	assign w29558 = w29460 ^ w29461;
	assign w29457 = w29453 ^ w29458;
	assign w29557 = w29456 ^ w29457;
	assign w29491 = w29521 & w29547;
	assign w29556 = w29481 ^ w29455;
	assign w29450 = ~w29454;
	assign w29452 = w29453 ^ w29491;
	assign w45670 = ~w29556;
	assign w43440 = w45317 ^ w45670;
	assign w45671 = ~w29557;
	assign w43447 = w45310 ^ w45671;
	assign w45672 = ~w29558;
	assign w43467 = w45311 ^ w45672;
	assign w29448 = w29452 ^ w44607;
	assign w29451 = w29490 ^ w29448;
	assign w29555 = w29450 ^ w29451;
	assign w45677 = ~w29555;
	assign w29446 = ~w29449;
	assign w29447 = w29471 ^ w29448;
	assign w50315 = w29446 ^ w29447;
	assign w43435 = w50311 ^ w50315;
	assign w29444 = w29500 ^ w29501;
	assign w29445 = w29503 ^ w29476;
	assign w50316 = w29444 ^ w29445;
	assign w43224 = w43417 ^ w50316;
	assign w43489 = w43224 ^ w43225;
	assign w43186 = w50316 ^ w50315;
	assign w45945 = ~w9484;
	assign w9279 = w45945 ^ w50060;
	assign w9552 = w9279 ^ w9280;
	assign w9316 = w45945 ^ w45339;
	assign w49944 = w9552 ^ w9549;
	assign w46713 = w49944 ^ w1209;
	assign w29731 = w46715 ^ w46713;
	assign w29733 = w46714 ^ w29731;
	assign w29808 = w29738 ^ w29733;
	assign w29806 = w46711 ^ w29733;
	assign w29802 = w29821 & w29806;
	assign w29809 = w46710 ^ w29733;
	assign w29736 = w29802 ^ w29732;
	assign w9403 = w45945 ^ w50058;
	assign w49945 = w9402 ^ w9403;
	assign w46712 = w49945 ^ w1210;
	assign w29822 = w46714 ^ w46712;
	assign w29807 = w29732 ^ w29822;
	assign w29798 = w29822 & w29807;
	assign w29734 = w46712 ^ w46710;
	assign w29693 = w29734 ^ w46711;
	assign w29817 = w46716 ^ w29693;
	assign w29803 = w46716 & w29817;
	assign w29694 = w29734 ^ w29732;
	assign w29810 = w29731 ^ w29694;
	assign w29797 = w29819 & w29810;
	assign w49924 = w9316 ^ w9317;
	assign w46733 = w49924 ^ w1189;
	assign w15749 = w46733 ^ w46738;
	assign w15751 = w46733 ^ w46739;
	assign w15662 = w46735 ^ w46733;
	assign w15745 = w15662 ^ w15668;
	assign w15743 = w15678 ^ w15745;
	assign w15730 = w15745 & w15738;
	assign w15624 = w15664 ^ w15662;
	assign w15740 = w15661 ^ w15624;
	assign w15727 = w15749 & w15740;
	assign w44025 = w15727 ^ w15733;
	assign w15677 = w44025 ^ w15662;
	assign w44026 = w15727 ^ w15730;
	assign w15750 = w46736 ^ w46733;
	assign w15729 = w15750 & w15739;
	assign w15746 = w15750 ^ w15678;
	assign w15665 = w15729 ^ w15663;
	assign w15742 = w15661 ^ w15750;
	assign w15735 = w15742 & w15746;
	assign w15667 = w15735 ^ w15664;
	assign w15671 = w15667 ^ w15665;
	assign w15676 = w46733 ^ w15671;
	assign w15741 = w46740 ^ w15742;
	assign w15734 = w15743 & w15741;
	assign w15639 = w15671 ^ w44025;
	assign w15682 = w46735 ^ w15639;
	assign w29820 = w46712 ^ w46709;
	assign w29799 = w29820 & w29809;
	assign w29816 = w29820 ^ w29748;
	assign w29735 = w29799 ^ w29733;
	assign w29707 = w29798 ^ w29799;
	assign w29812 = w29731 ^ w29820;
	assign w29811 = w46716 ^ w29812;
	assign w29805 = w29812 & w29816;
	assign w29737 = w29805 ^ w29734;
	assign w29741 = w29737 ^ w29735;
	assign w29746 = w46709 ^ w29741;
	assign w29800 = w29815 & w29808;
	assign w44615 = w29797 ^ w29803;
	assign w29709 = w29741 ^ w44615;
	assign w29752 = w46711 ^ w29709;
	assign w44616 = w29797 ^ w29800;
	assign w29750 = w29798 ^ w44616;
	assign w29710 = w29736 ^ w44616;
	assign w29794 = w29710 ^ w29735;
	assign w29706 = w29801 ^ w29750;
	assign w29788 = w46715 ^ w29706;
	assign w29804 = w29813 & w29811;
	assign w15737 = w15662 ^ w15752;
	assign w15728 = w15752 & w15737;
	assign w15637 = w15728 ^ w15729;
	assign w15680 = w15728 ^ w44026;
	assign w15636 = w15731 ^ w15680;
	assign w15684 = w15637 ^ w15638;
	assign w15718 = w46739 ^ w15636;
	assign w15685 = w15728 ^ w15734;
	assign w15723 = w15685 ^ w15677;
	assign w15726 = w15685 ^ w15676;
	assign w15732 = w15751 & w15736;
	assign w15666 = w15732 ^ w15662;
	assign w15640 = w15666 ^ w44026;
	assign w15724 = w15640 ^ w15665;
	assign w15683 = w15684 ^ w15666;
	assign w15725 = w15731 ^ w15683;
	assign w15722 = w15726 & w15725;
	assign w15717 = w15722 ^ w15682;
	assign w15716 = w15717 & w15718;
	assign w15715 = w15716 ^ w15724;
	assign w15634 = w15716 ^ w15733;
	assign w15629 = w15634 ^ w15730;
	assign w15701 = w15715 & w46740;
	assign w15721 = w15722 ^ w15724;
	assign w15720 = w15723 & w15721;
	assign w15719 = w15720 ^ w15682;
	assign w15631 = w15720 ^ w15732;
	assign w15627 = w15631 ^ w15667;
	assign w15689 = w15719 & w15745;
	assign w15630 = w46733 ^ w15627;
	assign w15707 = w15629 ^ w15630;
	assign w15688 = w15707 & w15750;
	assign w15628 = w15720 ^ w15676;
	assign w15698 = w15719 & w15738;
	assign w15635 = w15716 ^ w15680;
	assign w15692 = w15715 & w15747;
	assign w15626 = w46735 ^ w15627;
	assign w15714 = w15722 ^ w15716;
	assign w15713 = w15724 & w15714;
	assign w44029 = w15713 ^ w15731;
	assign w15672 = w46739 ^ w44029;
	assign w15712 = w15672 ^ w15635;
	assign w15693 = w15712 & w15743;
	assign w15705 = w44029 ^ w15683;
	assign w15694 = w15705 & w15746;
	assign w15703 = w15705 & w15742;
	assign w44028 = w15701 ^ w15703;
	assign w15702 = w15712 & w15741;
	assign w15697 = w15707 & w15739;
	assign w29747 = w44615 ^ w29732;
	assign w29708 = w46713 ^ w46714;
	assign w29754 = w29707 ^ w29708;
	assign w29753 = w29754 ^ w29736;
	assign w29795 = w29801 ^ w29753;
	assign w29755 = w29798 ^ w29804;
	assign w29796 = w29755 ^ w29746;
	assign w29792 = w29796 & w29795;
	assign w29787 = w29792 ^ w29752;
	assign w29786 = w29787 & w29788;
	assign w29785 = w29786 ^ w29794;
	assign w29762 = w29785 & w29817;
	assign w29771 = w29785 & w46716;
	assign w29704 = w29786 ^ w29803;
	assign w29784 = w29792 ^ w29786;
	assign w29783 = w29794 & w29784;
	assign w29705 = w29786 ^ w29750;
	assign w44619 = w29783 ^ w29801;
	assign w29742 = w46715 ^ w44619;
	assign w29775 = w44619 ^ w29753;
	assign w29764 = w29775 & w29816;
	assign w29773 = w29775 & w29812;
	assign w44618 = w29771 ^ w29773;
	assign w29782 = w29742 ^ w29705;
	assign w29772 = w29782 & w29811;
	assign w29763 = w29782 & w29813;
	assign w29699 = w29704 ^ w29800;
	assign w29791 = w29792 ^ w29794;
	assign w29781 = w29783 ^ w29791;
	assign w29793 = w29755 ^ w29747;
	assign w29790 = w29793 & w29791;
	assign w29789 = w29790 ^ w29752;
	assign w29759 = w29789 & w29815;
	assign w29698 = w29790 ^ w29746;
	assign w29701 = w29790 ^ w29802;
	assign w29768 = w29789 & w29808;
	assign w29697 = w29701 ^ w29737;
	assign w29780 = w29789 & w29781;
	assign w29745 = w29780 ^ w29755;
	assign w29779 = w29745 ^ w29747;
	assign w29760 = w29779 & w29814;
	assign w29769 = w29779 & w29818;
	assign w29712 = w29768 ^ w29769;
	assign w29703 = w29780 ^ w29804;
	assign w29695 = w29742 ^ w29703;
	assign w29702 = w29732 ^ w29695;
	assign w29778 = w29699 ^ w29702;
	assign w29765 = w29778 & w29810;
	assign w29730 = w29768 ^ w29760;
	assign w29776 = w29745 ^ w29698;
	assign w29761 = w29776 & w29821;
	assign w29743 = w29761 ^ w29765;
	assign w29721 = ~w29743;
	assign w29720 = w29721 ^ w29759;
	assign w29756 = w29778 & w29819;
	assign w29700 = w46709 ^ w29697;
	assign w29777 = w29699 ^ w29700;
	assign w29767 = w29777 & w29809;
	assign w29696 = w46711 ^ w29697;
	assign w29774 = w29695 ^ w29696;
	assign w29757 = w29774 & w29822;
	assign w29766 = w29774 & w29807;
	assign w29727 = w29766 ^ w29769;
	assign w29724 = ~w29727;
	assign w29758 = w29777 & w29820;
	assign w43582 = w29757 ^ w29758;
	assign w29726 = w29730 ^ w43582;
	assign w29729 = w44618 ^ w29726;
	assign w29725 = w29721 ^ w29726;
	assign w29825 = w29724 ^ w29725;
	assign w29716 = w29720 ^ w44618;
	assign w29719 = w29758 ^ w29716;
	assign w29770 = w29776 & w29806;
	assign w29728 = w29770 ^ w29761;
	assign w29826 = w29728 ^ w29729;
	assign w44617 = w29769 ^ w29770;
	assign w29751 = w29766 ^ w44617;
	assign w29717 = w29762 ^ w29751;
	assign w29714 = ~w29717;
	assign w29711 = w29767 ^ w29751;
	assign w29723 = w29766 ^ w29767;
	assign w29722 = w29767 ^ w29756;
	assign w29718 = ~w29722;
	assign w29823 = w29718 ^ w29719;
	assign w15711 = w15713 ^ w15721;
	assign w15710 = w15719 & w15711;
	assign w15675 = w15710 ^ w15685;
	assign w15706 = w15675 ^ w15628;
	assign w15709 = w15675 ^ w15677;
	assign w15690 = w15709 & w15744;
	assign w15660 = w15698 ^ w15690;
	assign w15699 = w15709 & w15748;
	assign w15642 = w15698 ^ w15699;
	assign w15633 = w15710 ^ w15734;
	assign w15700 = w15706 & w15736;
	assign w44027 = w15699 ^ w15700;
	assign w15625 = w15672 ^ w15633;
	assign w15632 = w15662 ^ w15625;
	assign w15708 = w15629 ^ w15632;
	assign w15704 = w15625 ^ w15626;
	assign w15696 = w15704 & w15737;
	assign w15681 = w15696 ^ w44027;
	assign w15687 = w15704 & w15752;
	assign w15657 = w15696 ^ w15699;
	assign w15641 = w15697 ^ w15681;
	assign w15654 = ~w15657;
	assign w15686 = w15708 & w15749;
	assign w43542 = w15687 ^ w15688;
	assign w15656 = w15660 ^ w43542;
	assign w15695 = w15708 & w15740;
	assign w15647 = w15692 ^ w15681;
	assign w15644 = ~w15647;
	assign w15653 = w15696 ^ w15697;
	assign w15669 = w15693 ^ w43542;
	assign w15670 = w15694 ^ w15669;
	assign w15674 = w15702 ^ w15670;
	assign w15679 = w15703 ^ w15674;
	assign w15659 = w44028 ^ w15656;
	assign w15652 = w15697 ^ w15686;
	assign w15648 = ~w15652;
	assign w15754 = w15679 ^ w15653;
	assign w50305 = ~w15754;
	assign w15643 = w15701 ^ w15674;
	assign w50304 = w44027 ^ w15679;
	assign w43223 = ~w50304;
	assign w43412 = w50317 ^ w43223;
	assign w50306 = w15670 ^ w15641;
	assign w43429 = w50306 ^ w50318;
	assign w43228 = w43467 ^ w43429;
	assign w29739 = w29763 ^ w43582;
	assign w29740 = w29764 ^ w29739;
	assign w50265 = w29740 ^ w29711;
	assign w43423 = w50260 ^ w50265;
	assign w43431 = w50249 ^ w50265;
	assign w43416 = w43464 ^ w43431;
	assign w43365 = w43474 ^ w43423;
	assign w50133 = w50249 ^ w43365;
	assign w43327 = ~w43431;
	assign w43347 = w43464 ^ w43423;
	assign w50142 = w45319 ^ w43347;
	assign w46588 = w50142 ^ w1333;
	assign w43326 = w43327 ^ w50251;
	assign w43173 = w43431 ^ w50247;
	assign w46597 = w50133 ^ w1324;
	assign w29744 = w29772 ^ w29740;
	assign w29713 = w29771 ^ w29744;
	assign w29715 = w29739 ^ w29716;
	assign w50261 = w29714 ^ w29715;
	assign w43466 = w50246 ^ w50261;
	assign w43328 = ~w43466;
	assign w43397 = w43328 ^ w45227;
	assign w50128 = w43397 ^ w43398;
	assign w43360 = w43466 ^ w43465;
	assign w50136 = w50250 ^ w43360;
	assign w46594 = w50136 ^ w1327;
	assign w46602 = w50128 ^ w1319;
	assign w32901 = w46597 ^ w46602;
	assign w29749 = w29773 ^ w29744;
	assign w29824 = w29749 ^ w29723;
	assign w50264 = ~w29824;
	assign w50263 = w44617 ^ w29749;
	assign w43468 = w45589 ^ w50264;
	assign w43475 = w50259 ^ w50263;
	assign w43368 = w43370 ^ w43475;
	assign w43366 = w43476 ^ w43468;
	assign w50132 = w45325 ^ w43366;
	assign w46598 = w50132 ^ w1323;
	assign w43350 = w43474 ^ w29824;
	assign w50140 = w43350 ^ w43351;
	assign w46590 = w50140 ^ w1331;
	assign w43340 = w43476 ^ w43475;
	assign w50147 = w45588 ^ w43340;
	assign w46583 = w50147 ^ w1338;
	assign w43337 = w43468 ^ w43424;
	assign w50149 = w50260 ^ w43337;
	assign w43293 = w50263 ^ w11331;
	assign w43275 = w43468 ^ w45324;
	assign w43256 = w29824 ^ w50255;
	assign w43210 = w43425 ^ w50263;
	assign w43495 = w43210 ^ w43211;
	assign w50138 = w43495 ^ w43479;
	assign w46592 = w50138 ^ w1329;
	assign w14948 = w46594 ^ w46592;
	assign w46581 = w50149 ^ w1340;
	assign w29330 = w46583 ^ w46581;
	assign w14860 = w46592 ^ w46590;
	assign w50262 = w29712 ^ w29713;
	assign w43478 = w50258 ^ w50262;
	assign w50129 = w43493 ^ w43478;
	assign w46601 = w50129 ^ w1320;
	assign w32790 = w46601 ^ w46602;
	assign w43358 = w43359 ^ w50262;
	assign w50137 = w43357 ^ w43358;
	assign w43343 = w43479 ^ w43478;
	assign w43341 = ~w43343;
	assign w43325 = w43478 ^ w43328;
	assign w50121 = w43325 ^ w43326;
	assign w46609 = w50121 ^ w1312;
	assign w43174 = w50262 ^ w50252;
	assign w43510 = w43173 ^ w43174;
	assign w50122 = w43510 ^ w43475;
	assign w46608 = w50122 ^ w1313;
	assign w46593 = w50137 ^ w1328;
	assign w14834 = w46593 ^ w46594;
	assign w45678 = ~w29823;
	assign w43471 = w45588 ^ w45678;
	assign w43367 = w43479 ^ w43471;
	assign w50131 = w45324 ^ w43367;
	assign w46599 = w50131 ^ w1322;
	assign w32814 = w46599 ^ w46597;
	assign w43352 = w43476 ^ w45678;
	assign w50139 = w43352 ^ w43353;
	assign w46591 = w50139 ^ w1330;
	assign w43338 = w43474 ^ w43471;
	assign w50148 = w45589 ^ w43338;
	assign w46582 = w50148 ^ w1339;
	assign w29336 = w46588 ^ w46582;
	assign w29416 = w46583 ^ w29336;
	assign w43294 = w43471 ^ w50248;
	assign w43292 = ~w43294;
	assign w50123 = w43292 ^ w43293;
	assign w46607 = w50123 ^ w1314;
	assign w43276 = w45678 ^ w11332;
	assign w43274 = w43275 ^ w43276;
	assign w50124 = ~w43274;
	assign w46606 = w50124 ^ w1315;
	assign w29413 = w29330 ^ w29336;
	assign w14994 = w46608 ^ w46606;
	assign w14953 = w14994 ^ w46607;
	assign w14819 = w14860 ^ w46591;
	assign w45679 = ~w29825;
	assign w43486 = w45318 ^ w45679;
	assign w43362 = w43486 ^ w43464;
	assign w43361 = w43362 ^ w43363;
	assign w50135 = ~w43361;
	assign w43356 = w43327 ^ w45679;
	assign w43345 = w45679 ^ w26475;
	assign w50144 = w43344 ^ w43345;
	assign w46586 = w50144 ^ w1335;
	assign w29417 = w46581 ^ w46586;
	assign w43339 = w43486 ^ w43463;
	assign w50120 = w50261 ^ w43339;
	assign w46610 = w50120 ^ w1311;
	assign w14968 = w46609 ^ w46610;
	assign w15082 = w46610 ^ w46608;
	assign w46595 = w50135 ^ w1326;
	assign w14857 = w46595 ^ w46593;
	assign w14859 = w46594 ^ w14857;
	assign w14874 = w46595 ^ w46594;
	assign w14932 = w46591 ^ w14859;
	assign w14935 = w46590 ^ w14859;
	assign w45680 = ~w29826;
	assign w43487 = w45319 ^ w45680;
	assign w50118 = w45680 ^ w43416;
	assign w46612 = w50118 ^ w1309;
	assign w15077 = w46612 ^ w14953;
	assign w14998 = w46612 ^ w46606;
	assign w15078 = w46607 ^ w14998;
	assign w15063 = w46612 & w15077;
	assign w43364 = w43487 ^ w43425;
	assign w50134 = w45228 ^ w43364;
	assign w46596 = w50134 ^ w1325;
	assign w14864 = w46596 ^ w46590;
	assign w14944 = w46591 ^ w14864;
	assign w14934 = w14864 ^ w14859;
	assign w14943 = w46596 ^ w14819;
	assign w14940 = w46595 ^ w14944;
	assign w14927 = w14944 & w14940;
	assign w14929 = w46596 & w14943;
	assign w43355 = w43487 ^ w43465;
	assign w43354 = w43355 ^ w43356;
	assign w50119 = ~w43354;
	assign w43239 = w43487 ^ w43424;
	assign w50126 = w45582 ^ w43239;
	assign w46604 = w50126 ^ w1317;
	assign w32820 = w46604 ^ w46598;
	assign w32897 = w32814 ^ w32820;
	assign w32900 = w46599 ^ w32820;
	assign w43216 = w43423 ^ w45680;
	assign w43492 = w43216 ^ w43217;
	assign w50143 = w43492 ^ w43465;
	assign w46587 = w50143 ^ w1334;
	assign w29346 = w46587 ^ w46586;
	assign w29412 = w46587 ^ w29416;
	assign w29399 = w29416 & w29412;
	assign w29411 = w29346 ^ w29413;
	assign w29419 = w46581 ^ w46587;
	assign w46611 = w50119 ^ w1310;
	assign w14991 = w46611 ^ w46609;
	assign w15074 = w46611 ^ w15078;
	assign w15061 = w15078 & w15074;
	assign w15008 = w46611 ^ w46610;
	assign w14993 = w46610 ^ w14991;
	assign w15069 = w46606 ^ w14993;
	assign w15066 = w46607 ^ w14993;
	assign w15068 = w14998 ^ w14993;
	assign w50303 = w15642 ^ w15643;
	assign w43443 = w50303 ^ w50316;
	assign w43414 = w43443 ^ w43434;
	assign w15691 = w15706 & w15751;
	assign w15658 = w15700 ^ w15691;
	assign w15756 = w15658 ^ w15659;
	assign w45323 = ~w15756;
	assign w43183 = w43429 ^ w45323;
	assign w15673 = w15691 ^ w15695;
	assign w15651 = ~w15673;
	assign w15650 = w15651 ^ w15689;
	assign w15646 = w15650 ^ w44028;
	assign w15655 = w15651 ^ w15656;
	assign w15649 = w15688 ^ w15646;
	assign w15753 = w15648 ^ w15649;
	assign w15755 = w15654 ^ w15655;
	assign w15645 = w15669 ^ w15646;
	assign w50302 = w15644 ^ w15645;
	assign w43185 = w43429 ^ w50302;
	assign w43505 = w43185 ^ w43186;
	assign w45322 = ~w15755;
	assign w43226 = w43435 ^ w45322;
	assign w45329 = ~w15753;
	assign w43452 = w45329 ^ w45677;
	assign w43410 = w43452 ^ w43440;
	assign w43396 = w15754 ^ w45329;
	assign w43386 = w43452 ^ w50313;
	assign w45946 = ~w9482;
	assign w9380 = w45946 ^ w50066;
	assign w9384 = w45946 ^ w45336;
	assign w9382 = w9383 ^ w9384;
	assign w49958 = ~w9382;
	assign w46699 = w49958 ^ w1159;
	assign w33030 = w46699 ^ w33034;
	assign w33017 = w33034 & w33030;
	assign w33037 = w46693 ^ w46699;
	assign w32964 = w46699 ^ w46698;
	assign w33029 = w32964 ^ w33031;
	assign w49960 = w9379 ^ w9380;
	assign w46697 = w49960 ^ w1161;
	assign w32924 = w46697 ^ w46698;
	assign w32947 = w46699 ^ w46697;
	assign w9377 = w45946 ^ w50067;
	assign w49961 = w9376 ^ w9377;
	assign w46696 = w49961 ^ w1162;
	assign w33038 = w46698 ^ w46696;
	assign w33036 = w46696 ^ w46693;
	assign w33032 = w33036 ^ w32964;
	assign w33023 = w32948 ^ w33038;
	assign w33028 = w32947 ^ w33036;
	assign w33027 = w46700 ^ w33028;
	assign w33020 = w33029 & w33027;
	assign w33021 = w33028 & w33032;
	assign w32949 = w46698 ^ w32947;
	assign w33022 = w46695 ^ w32949;
	assign w33018 = w33037 & w33022;
	assign w32952 = w33018 ^ w32948;
	assign w33024 = w32954 ^ w32949;
	assign w33016 = w33031 & w33024;
	assign w33025 = w46694 ^ w32949;
	assign w33015 = w33036 & w33025;
	assign w32951 = w33015 ^ w32949;
	assign w32950 = w46696 ^ w46694;
	assign w32953 = w33021 ^ w32950;
	assign w32910 = w32950 ^ w32948;
	assign w32909 = w32950 ^ w46695;
	assign w33026 = w32947 ^ w32910;
	assign w33013 = w33035 & w33026;
	assign w33033 = w46700 ^ w32909;
	assign w33019 = w46700 & w33033;
	assign w44749 = w33013 ^ w33016;
	assign w32926 = w32952 ^ w44749;
	assign w33010 = w32926 ^ w32951;
	assign w44752 = w33013 ^ w33019;
	assign w32963 = w44752 ^ w32948;
	assign w32957 = w32953 ^ w32951;
	assign w32925 = w32957 ^ w44752;
	assign w32962 = w46693 ^ w32957;
	assign w32968 = w46695 ^ w32925;
	assign w33014 = w33038 & w33023;
	assign w32966 = w33014 ^ w44749;
	assign w32923 = w33014 ^ w33015;
	assign w32970 = w32923 ^ w32924;
	assign w32969 = w32970 ^ w32952;
	assign w33011 = w33017 ^ w32969;
	assign w32922 = w33017 ^ w32966;
	assign w33004 = w46699 ^ w32922;
	assign w32971 = w33014 ^ w33020;
	assign w33009 = w32971 ^ w32963;
	assign w33012 = w32971 ^ w32962;
	assign w33008 = w33012 & w33011;
	assign w33007 = w33008 ^ w33010;
	assign w33003 = w33008 ^ w32968;
	assign w33002 = w33003 & w33004;
	assign w32920 = w33002 ^ w33019;
	assign w32915 = w32920 ^ w33016;
	assign w33001 = w33002 ^ w33010;
	assign w32987 = w33001 & w46700;
	assign w32921 = w33002 ^ w32966;
	assign w33000 = w33008 ^ w33002;
	assign w32999 = w33010 & w33000;
	assign w33006 = w33009 & w33007;
	assign w32917 = w33006 ^ w33018;
	assign w32913 = w32917 ^ w32953;
	assign w32912 = w46695 ^ w32913;
	assign w32914 = w33006 ^ w32962;
	assign w33005 = w33006 ^ w32968;
	assign w32984 = w33005 & w33024;
	assign w32978 = w33001 & w33033;
	assign w32997 = w32999 ^ w33007;
	assign w32996 = w33005 & w32997;
	assign w32961 = w32996 ^ w32971;
	assign w32919 = w32996 ^ w33020;
	assign w32992 = w32961 ^ w32914;
	assign w32995 = w32961 ^ w32963;
	assign w32985 = w32995 & w33034;
	assign w32928 = w32984 ^ w32985;
	assign w32986 = w32992 & w33022;
	assign w44751 = w32999 ^ w33017;
	assign w32991 = w44751 ^ w32969;
	assign w32980 = w32991 & w33032;
	assign w32958 = w46699 ^ w44751;
	assign w32998 = w32958 ^ w32921;
	assign w32911 = w32958 ^ w32919;
	assign w32918 = w32948 ^ w32911;
	assign w32994 = w32915 ^ w32918;
	assign w32990 = w32911 ^ w32912;
	assign w32973 = w32990 & w33038;
	assign w32981 = w32994 & w33026;
	assign w32982 = w32990 & w33023;
	assign w32943 = w32982 ^ w32985;
	assign w32940 = ~w32943;
	assign w32972 = w32994 & w33035;
	assign w32979 = w32998 & w33029;
	assign w44753 = w32985 ^ w32986;
	assign w32967 = w32982 ^ w44753;
	assign w32933 = w32978 ^ w32967;
	assign w32930 = ~w32933;
	assign w32916 = w46693 ^ w32913;
	assign w32993 = w32915 ^ w32916;
	assign w32983 = w32993 & w33025;
	assign w32939 = w32982 ^ w32983;
	assign w32938 = w32983 ^ w32972;
	assign w32934 = ~w32938;
	assign w32927 = w32983 ^ w32967;
	assign w32989 = w32991 & w33028;
	assign w44754 = w32987 ^ w32989;
	assign w32988 = w32998 & w33027;
	assign w32977 = w32992 & w33037;
	assign w32944 = w32986 ^ w32977;
	assign w32959 = w32977 ^ w32981;
	assign w32937 = ~w32959;
	assign w32976 = w32995 & w33030;
	assign w32946 = w32984 ^ w32976;
	assign w32975 = w33005 & w33031;
	assign w32936 = w32937 ^ w32975;
	assign w32932 = w32936 ^ w44754;
	assign w32974 = w32993 & w33036;
	assign w32935 = w32974 ^ w32932;
	assign w33039 = w32934 ^ w32935;
	assign w44750 = w32973 ^ w32974;
	assign w32955 = w32979 ^ w44750;
	assign w32931 = w32955 ^ w32932;
	assign w50307 = w32930 ^ w32931;
	assign w43227 = w45671 ^ w50307;
	assign w50216 = w43226 ^ w43227;
	assign w46514 = w50216 ^ w1216;
	assign w43457 = w50302 ^ w50307;
	assign w43402 = w43457 ^ w43443;
	assign w43400 = ~w43402;
	assign w43390 = w43457 ^ w50315;
	assign w43378 = w43457 ^ w43447;
	assign w50240 = w50311 ^ w43378;
	assign w46490 = w50240 ^ w1240;
	assign w32942 = w32946 ^ w44750;
	assign w32941 = w32937 ^ w32942;
	assign w33041 = w32940 ^ w32941;
	assign w32945 = w44754 ^ w32942;
	assign w33042 = w32944 ^ w32945;
	assign w32956 = w32980 ^ w32955;
	assign w50310 = w32956 ^ w32927;
	assign w32960 = w32988 ^ w32956;
	assign w32965 = w32989 ^ w32960;
	assign w33040 = w32965 ^ w32939;
	assign w32929 = w32987 ^ w32960;
	assign w50308 = w32928 ^ w32929;
	assign w50309 = w44753 ^ w32965;
	assign w43418 = w50306 ^ w50310;
	assign w43432 = w50310 ^ w50314;
	assign w43437 = w50308 ^ w50312;
	assign w50217 = w43505 ^ w43437;
	assign w46513 = w50217 ^ w1217;
	assign w14432 = w46513 ^ w46514;
	assign w43483 = w50304 ^ w50309;
	assign w50242 = w43489 ^ w43483;
	assign w46488 = w50242 ^ w45169;
	assign w43415 = w43429 ^ w50309;
	assign w50218 = w43414 ^ w43415;
	assign w46512 = w50218 ^ w1218;
	assign w43409 = w50310 ^ w15754;
	assign w43407 = w43467 ^ w43418;
	assign w50222 = w45323 ^ w43407;
	assign w46508 = w50222 ^ w1222;
	assign w43399 = w43483 ^ w43452;
	assign w50227 = w45316 ^ w43399;
	assign w46503 = w50227 ^ w1227;
	assign w43388 = w43483 ^ w43437;
	assign w43389 = w43432 ^ w50317;
	assign w50234 = w43388 ^ w43389;
	assign w46496 = w50234 ^ w1234;
	assign w43383 = w43418 ^ w50318;
	assign w43376 = w43437 ^ w43435;
	assign w43371 = w43440 ^ w43418;
	assign w50245 = w50314 ^ w43371;
	assign w46485 = w50245 ^ w1244;
	assign w29149 = w46485 ^ w46490;
	assign w29150 = w46488 ^ w46485;
	assign w43222 = w50308 ^ w43223;
	assign w43171 = w43432 ^ w50311;
	assign w43172 = w50308 ^ w50307;
	assign w43511 = w43171 ^ w43172;
	assign w50233 = w43511 ^ w43443;
	assign w46497 = w50233 ^ w1233;
	assign w43169 = w43432 ^ w45671;
	assign w29152 = w46490 ^ w46488;
	assign w45762 = ~w33042;
	assign w43480 = w45323 ^ w45762;
	assign w43405 = w43480 ^ w43447;
	assign w43392 = w43480 ^ w43432;
	assign w50230 = w45672 ^ w43392;
	assign w46500 = w50230 ^ w1230;
	assign w43382 = w43480 ^ w43417;
	assign w50238 = w45311 ^ w43382;
	assign w50214 = w45762 ^ w43228;
	assign w46516 = w50214 ^ w1214;
	assign w43170 = w45311 ^ w45762;
	assign w43512 = w43169 ^ w43170;
	assign w46492 = w50238 ^ w1238;
	assign w45767 = ~w33039;
	assign w43442 = w45767 ^ w45316;
	assign w43413 = ~w43442;
	assign w43411 = w43413 ^ w45677;
	assign w50219 = w43411 ^ w43412;
	assign w46511 = w50219 ^ w1219;
	assign w43395 = w43440 ^ w45767;
	assign w43394 = w43395 ^ w43396;
	assign w50228 = ~w43394;
	assign w46502 = w50228 ^ w1228;
	assign w32686 = w46508 ^ w46502;
	assign w32766 = w46503 ^ w32686;
	assign w43387 = w45767 ^ w50309;
	assign w50235 = w43386 ^ w43387;
	assign w46495 = w50235 ^ w1235;
	assign w43374 = w43442 ^ w43434;
	assign w50243 = w45329 ^ w43374;
	assign w46487 = w50243 ^ w1242;
	assign w29062 = w46487 ^ w46485;
	assign w29137 = w29062 ^ w29152;
	assign w29128 = w29152 & w29137;
	assign w45768 = ~w33040;
	assign w43482 = w50305 ^ w45768;
	assign w50220 = w45768 ^ w43410;
	assign w46510 = w50220 ^ w1220;
	assign w14462 = w46516 ^ w46510;
	assign w14542 = w46511 ^ w14462;
	assign w14458 = w46512 ^ w46510;
	assign w14417 = w14458 ^ w46511;
	assign w14541 = w46516 ^ w14417;
	assign w43393 = w43482 ^ w43417;
	assign w50229 = w50306 ^ w43393;
	assign w46501 = w50229 ^ w1229;
	assign w43385 = w43482 ^ w43442;
	assign w50236 = w45670 ^ w43385;
	assign w46494 = w50236 ^ w1236;
	assign w14328 = w46500 ^ w46494;
	assign w14408 = w46495 ^ w14328;
	assign w14324 = w46496 ^ w46494;
	assign w43384 = w45317 ^ w45768;
	assign w50237 = w43383 ^ w43384;
	assign w46493 = w50237 ^ w1237;
	assign w14322 = w46495 ^ w46493;
	assign w14410 = w46496 ^ w46493;
	assign w14405 = w14322 ^ w14328;
	assign w14284 = w14324 ^ w14322;
	assign w43372 = w43482 ^ w45677;
	assign w50244 = w43372 ^ w43373;
	assign w46486 = w50244 ^ w1243;
	assign w29068 = w46492 ^ w46486;
	assign w29148 = w46487 ^ w29068;
	assign w14283 = w14324 ^ w46495;
	assign w14407 = w46500 ^ w14283;
	assign w14393 = w46500 & w14407;
	assign w14527 = w46516 & w14541;
	assign w29145 = w29062 ^ w29068;
	assign w29064 = w46488 ^ w46486;
	assign w29024 = w29064 ^ w29062;
	assign w29023 = w29064 ^ w46487;
	assign w29147 = w46492 ^ w29023;
	assign w29133 = w46492 & w29147;
	assign w32680 = w46503 ^ w46501;
	assign w32763 = w32680 ^ w32686;
	assign w45769 = ~w33041;
	assign w43472 = w45322 ^ w45769;
	assign w50231 = w43512 ^ w43472;
	assign w46499 = w50231 ^ w1231;
	assign w14321 = w46499 ^ w46497;
	assign w14402 = w14321 ^ w14410;
	assign w14401 = w46500 ^ w14402;
	assign w14411 = w46493 ^ w46499;
	assign w14404 = w46499 ^ w14408;
	assign w14391 = w14408 & w14404;
	assign w14400 = w14321 ^ w14284;
	assign w43403 = w43472 ^ w43435;
	assign w50224 = w50302 ^ w43403;
	assign w46506 = w50224 ^ w1224;
	assign w32767 = w46501 ^ w46506;
	assign w43391 = w45310 ^ w45769;
	assign w50232 = w43390 ^ w43391;
	assign w43381 = ~w43472;
	assign w43379 = w43381 ^ w43467;
	assign w43184 = w45672 ^ w45769;
	assign w43506 = w43183 ^ w43184;
	assign w50215 = w43506 ^ w43447;
	assign w46515 = w50215 ^ w1215;
	assign w14455 = w46515 ^ w46513;
	assign w14538 = w46515 ^ w14542;
	assign w14525 = w14542 & w14538;
	assign w14472 = w46515 ^ w46514;
	assign w14457 = w46514 ^ w14455;
	assign w14532 = w14462 ^ w14457;
	assign w14530 = w46511 ^ w14457;
	assign w46498 = w50232 ^ w1232;
	assign w14409 = w46493 ^ w46498;
	assign w14338 = w46499 ^ w46498;
	assign w14298 = w46497 ^ w46498;
	assign w14412 = w46498 ^ w46496;
	assign w14397 = w14322 ^ w14412;
	assign w14388 = w14412 & w14397;
	assign w14406 = w14410 ^ w14338;
	assign w14403 = w14338 ^ w14405;
	assign w14394 = w14403 & w14401;
	assign w14395 = w14402 & w14406;
	assign w14327 = w14395 ^ w14324;
	assign w14323 = w46498 ^ w14321;
	assign w14398 = w14328 ^ w14323;
	assign w14390 = w14405 & w14398;
	assign w14399 = w46494 ^ w14323;
	assign w14389 = w14410 & w14399;
	assign w14325 = w14389 ^ w14323;
	assign w14297 = w14388 ^ w14389;
	assign w14344 = w14297 ^ w14298;
	assign w14331 = w14327 ^ w14325;
	assign w14336 = w46493 ^ w14331;
	assign w14396 = w46495 ^ w14323;
	assign w14392 = w14411 & w14396;
	assign w14326 = w14392 ^ w14322;
	assign w14343 = w14344 ^ w14326;
	assign w14385 = w14391 ^ w14343;
	assign w14533 = w46510 ^ w14457;
	assign w14345 = w14388 ^ w14394;
	assign w14386 = w14345 ^ w14336;
	assign w14382 = w14386 & w14385;
	assign w14387 = w14409 & w14400;
	assign w43969 = w14387 ^ w14390;
	assign w14340 = w14388 ^ w43969;
	assign w14296 = w14391 ^ w14340;
	assign w43972 = w14387 ^ w14393;
	assign w14299 = w14331 ^ w43972;
	assign w14342 = w46495 ^ w14299;
	assign w14377 = w14382 ^ w14342;
	assign w14337 = w43972 ^ w14322;
	assign w14383 = w14345 ^ w14337;
	assign w14378 = w46499 ^ w14296;
	assign w14376 = w14377 & w14378;
	assign w14374 = w14382 ^ w14376;
	assign w14295 = w14376 ^ w14340;
	assign w14294 = w14376 ^ w14393;
	assign w14289 = w14294 ^ w14390;
	assign w14300 = w14326 ^ w43969;
	assign w14384 = w14300 ^ w14325;
	assign w14381 = w14382 ^ w14384;
	assign w14373 = w14384 & w14374;
	assign w14371 = w14373 ^ w14381;
	assign w14380 = w14383 & w14381;
	assign w14379 = w14380 ^ w14342;
	assign w14349 = w14379 & w14405;
	assign w14370 = w14379 & w14371;
	assign w14293 = w14370 ^ w14394;
	assign w14291 = w14380 ^ w14392;
	assign w14375 = w14376 ^ w14384;
	assign w14288 = w14380 ^ w14336;
	assign w14361 = w14375 & w46500;
	assign w14358 = w14379 & w14398;
	assign w14352 = w14375 & w14407;
	assign w43971 = w14373 ^ w14391;
	assign w14365 = w43971 ^ w14343;
	assign w14363 = w14365 & w14402;
	assign w14354 = w14365 & w14406;
	assign w14332 = w46499 ^ w43971;
	assign w14285 = w14332 ^ w14293;
	assign w14292 = w14322 ^ w14285;
	assign w14372 = w14332 ^ w14295;
	assign w14368 = w14289 ^ w14292;
	assign w14355 = w14368 & w14400;
	assign w14353 = w14372 & w14403;
	assign w14362 = w14372 & w14401;
	assign w14346 = w14368 & w14409;
	assign w43974 = w14361 ^ w14363;
	assign w14335 = w14370 ^ w14345;
	assign w14366 = w14335 ^ w14288;
	assign w14369 = w14335 ^ w14337;
	assign w14360 = w14366 & w14396;
	assign w14359 = w14369 & w14408;
	assign w14302 = w14358 ^ w14359;
	assign w14351 = w14366 & w14411;
	assign w14318 = w14360 ^ w14351;
	assign w14333 = w14351 ^ w14355;
	assign w14311 = ~w14333;
	assign w14310 = w14311 ^ w14349;
	assign w14306 = w14310 ^ w43974;
	assign w43973 = w14359 ^ w14360;
	assign w14287 = w14291 ^ w14327;
	assign w14290 = w46493 ^ w14287;
	assign w14367 = w14289 ^ w14290;
	assign w14348 = w14367 & w14410;
	assign w14309 = w14348 ^ w14306;
	assign w14286 = w46495 ^ w14287;
	assign w14364 = w14285 ^ w14286;
	assign w14356 = w14364 & w14397;
	assign w14341 = w14356 ^ w43973;
	assign w14307 = w14352 ^ w14341;
	assign w14317 = w14356 ^ w14359;
	assign w14314 = ~w14317;
	assign w14347 = w14364 & w14412;
	assign w14357 = w14367 & w14399;
	assign w14313 = w14356 ^ w14357;
	assign w14312 = w14357 ^ w14346;
	assign w14308 = ~w14312;
	assign w14413 = w14308 ^ w14309;
	assign w14301 = w14357 ^ w14341;
	assign w43970 = w14347 ^ w14348;
	assign w14329 = w14353 ^ w43970;
	assign w14330 = w14354 ^ w14329;
	assign w14334 = w14362 ^ w14330;
	assign w14339 = w14363 ^ w14334;
	assign w50460 = w43973 ^ w14339;
	assign w14303 = w14361 ^ w14334;
	assign w50461 = w14330 ^ w14301;
	assign w50459 = w14302 ^ w14303;
	assign w14414 = w14339 ^ w14313;
	assign w14350 = w14369 & w14404;
	assign w14320 = w14358 ^ w14350;
	assign w14316 = w14320 ^ w43970;
	assign w14319 = w43974 ^ w14316;
	assign w14416 = w14318 ^ w14319;
	assign w14304 = ~w14307;
	assign w14315 = w14311 ^ w14316;
	assign w14415 = w14314 ^ w14315;
	assign w50457 = ~w14415;
	assign w14305 = w14329 ^ w14306;
	assign w50458 = w14304 ^ w14305;
	assign w42876 = ~w50458;
	assign w42875 = w50459 ^ w42876;
	assign w45287 = ~w14413;
	assign w45288 = ~w14414;
	assign w45289 = ~w14416;
	assign w14546 = w46514 ^ w46512;
	assign w45947 = ~w9480;
	assign w9302 = w45947 ^ w45598;
	assign w9297 = w45947 ^ w50094;
	assign w50008 = w9296 ^ w9297;
	assign w9294 = w45947 ^ w50095;
	assign w50009 = w9293 ^ w9294;
	assign w46648 = w50009 ^ w1146;
	assign w23790 = w46648 ^ w46645;
	assign w46649 = w50008 ^ w1145;
	assign w23678 = w46649 ^ w46650;
	assign w23792 = w46650 ^ w46648;
	assign w23777 = w23702 ^ w23792;
	assign w23768 = w23792 & w23777;
	assign w23704 = w46648 ^ w46646;
	assign w23664 = w23704 ^ w23702;
	assign w23663 = w23704 ^ w46647;
	assign w23787 = w46652 ^ w23663;
	assign w23773 = w46652 & w23787;
	assign w50006 = w9301 ^ w9302;
	assign w46651 = w50006 ^ w1143;
	assign w23701 = w46651 ^ w46649;
	assign w23782 = w23701 ^ w23790;
	assign w23780 = w23701 ^ w23664;
	assign w23781 = w46652 ^ w23782;
	assign w23767 = w23789 & w23780;
	assign w44363 = w23767 ^ w23773;
	assign w23718 = w46651 ^ w46650;
	assign w23783 = w23718 ^ w23785;
	assign w23774 = w23783 & w23781;
	assign w23786 = w23790 ^ w23718;
	assign w23725 = w23768 ^ w23774;
	assign w23775 = w23782 & w23786;
	assign w23707 = w23775 ^ w23704;
	assign w23717 = w44363 ^ w23702;
	assign w23763 = w23725 ^ w23717;
	assign w23703 = w46650 ^ w23701;
	assign w23779 = w46646 ^ w23703;
	assign w23769 = w23790 & w23779;
	assign w23705 = w23769 ^ w23703;
	assign w23711 = w23707 ^ w23705;
	assign w23716 = w46645 ^ w23711;
	assign w23766 = w23725 ^ w23716;
	assign w23679 = w23711 ^ w44363;
	assign w23722 = w46647 ^ w23679;
	assign w23677 = w23768 ^ w23769;
	assign w23724 = w23677 ^ w23678;
	assign w23778 = w23708 ^ w23703;
	assign w23770 = w23785 & w23778;
	assign w44364 = w23767 ^ w23770;
	assign w23791 = w46645 ^ w46651;
	assign w23776 = w46647 ^ w23703;
	assign w23772 = w23791 & w23776;
	assign w23706 = w23772 ^ w23702;
	assign w23723 = w23724 ^ w23706;
	assign w23680 = w23706 ^ w44364;
	assign w23764 = w23680 ^ w23705;
	assign w23784 = w46651 ^ w23788;
	assign w23771 = w23788 & w23784;
	assign w23765 = w23771 ^ w23723;
	assign w23762 = w23766 & w23765;
	assign w23757 = w23762 ^ w23722;
	assign w23761 = w23762 ^ w23764;
	assign w23760 = w23763 & w23761;
	assign w23759 = w23760 ^ w23722;
	assign w23738 = w23759 & w23778;
	assign w23729 = w23759 & w23785;
	assign w23668 = w23760 ^ w23716;
	assign w23671 = w23760 ^ w23772;
	assign w23667 = w23671 ^ w23707;
	assign w23670 = w46645 ^ w23667;
	assign w23666 = w46647 ^ w23667;
	assign w23720 = w23768 ^ w44364;
	assign w23676 = w23771 ^ w23720;
	assign w23758 = w46651 ^ w23676;
	assign w23756 = w23757 & w23758;
	assign w23754 = w23762 ^ w23756;
	assign w23755 = w23756 ^ w23764;
	assign w23732 = w23755 & w23787;
	assign w23675 = w23756 ^ w23720;
	assign w23741 = w23755 & w46652;
	assign w23674 = w23756 ^ w23773;
	assign w23669 = w23674 ^ w23770;
	assign w23747 = w23669 ^ w23670;
	assign w23728 = w23747 & w23790;
	assign w23737 = w23747 & w23779;
	assign w23753 = w23764 & w23754;
	assign w23751 = w23753 ^ w23761;
	assign w23750 = w23759 & w23751;
	assign w23673 = w23750 ^ w23774;
	assign w44367 = w23753 ^ w23771;
	assign w23745 = w44367 ^ w23723;
	assign w23743 = w23745 & w23782;
	assign w23734 = w23745 & w23786;
	assign w44366 = w23741 ^ w23743;
	assign w23712 = w46651 ^ w44367;
	assign w23752 = w23712 ^ w23675;
	assign w23742 = w23752 & w23781;
	assign w23733 = w23752 & w23783;
	assign w23665 = w23712 ^ w23673;
	assign w23744 = w23665 ^ w23666;
	assign w23736 = w23744 & w23777;
	assign w23693 = w23736 ^ w23737;
	assign w23672 = w23702 ^ w23665;
	assign w23748 = w23669 ^ w23672;
	assign w23735 = w23748 & w23780;
	assign w23726 = w23748 & w23789;
	assign w23692 = w23737 ^ w23726;
	assign w23688 = ~w23692;
	assign w23727 = w23744 & w23792;
	assign w43564 = w23727 ^ w23728;
	assign w23709 = w23733 ^ w43564;
	assign w23710 = w23734 ^ w23709;
	assign w23714 = w23742 ^ w23710;
	assign w23683 = w23741 ^ w23714;
	assign w23719 = w23743 ^ w23714;
	assign w23794 = w23719 ^ w23693;
	assign w45510 = ~w23794;
	assign w43433 = w45321 ^ w45510;
	assign w23715 = w23750 ^ w23725;
	assign w23746 = w23715 ^ w23668;
	assign w23740 = w23746 & w23776;
	assign w23749 = w23715 ^ w23717;
	assign w23730 = w23749 & w23784;
	assign w23700 = w23738 ^ w23730;
	assign w23696 = w23700 ^ w43564;
	assign w23699 = w44366 ^ w23696;
	assign w23731 = w23746 & w23791;
	assign w23713 = w23731 ^ w23735;
	assign w23698 = w23740 ^ w23731;
	assign w23796 = w23698 ^ w23699;
	assign w23691 = ~w23713;
	assign w23690 = w23691 ^ w23729;
	assign w23686 = w23690 ^ w44366;
	assign w23689 = w23728 ^ w23686;
	assign w23685 = w23709 ^ w23686;
	assign w23793 = w23688 ^ w23689;
	assign w23695 = w23691 ^ w23696;
	assign w45512 = ~w23796;
	assign w43481 = w45315 ^ w45512;
	assign w45517 = ~w23793;
	assign w43444 = w45320 ^ w45517;
	assign w43272 = w43433 ^ w45517;
	assign w23739 = w23749 & w23788;
	assign w23682 = w23738 ^ w23739;
	assign w50299 = w23682 ^ w23683;
	assign w23697 = w23736 ^ w23739;
	assign w23694 = ~w23697;
	assign w43459 = w50295 ^ w50299;
	assign w23795 = w23694 ^ w23695;
	assign w44365 = w23739 ^ w23740;
	assign w50300 = w44365 ^ w23719;
	assign w43450 = w50296 ^ w50300;
	assign w43279 = w43444 ^ w50300;
	assign w43277 = ~w43279;
	assign w23721 = w23736 ^ w44365;
	assign w23681 = w23737 ^ w23721;
	assign w50301 = w23710 ^ w23681;
	assign w23687 = w23732 ^ w23721;
	assign w23684 = ~w23687;
	assign w43419 = w50297 ^ w50301;
	assign w43427 = w50286 ^ w50301;
	assign w43283 = w43481 ^ w43427;
	assign w43269 = w43419 ^ w45510;
	assign w43200 = w43427 ^ w50299;
	assign w43196 = ~w43427;
	assign w43194 = w43196 ^ w45512;
	assign w50298 = w23684 ^ w23685;
	assign w43469 = w50294 ^ w50298;
	assign w43282 = ~w43469;
	assign w43197 = w43196 ^ w50298;
	assign w45511 = ~w23795;
	assign w43473 = w45314 ^ w45511;
	assign w43280 = w43282 ^ w45511;
	assign w45948 = ~w9479;
	assign w9282 = w45948 ^ w50102;
	assign w9551 = w9282 ^ w9283;
	assign w9467 = w45948 ^ w45602;
	assign w9465 = w9466 ^ w9467;
	assign w50022 = ~w9465;
	assign w9462 = w45948 ^ w50111;
	assign w50024 = w9461 ^ w9462;
	assign w46633 = w50024 ^ w1097;
	assign w46635 = w50022 ^ w1095;
	assign w11105 = w46635 ^ w46633;
	assign w11188 = w46635 ^ w11192;
	assign w11175 = w11192 & w11188;
	assign w11082 = w46633 ^ w46634;
	assign w50025 = w9551 ^ w9495;
	assign w11195 = w46629 ^ w46635;
	assign w46632 = w50025 ^ w1098;
	assign w11196 = w46634 ^ w46632;
	assign w11194 = w46632 ^ w46629;
	assign w11108 = w46632 ^ w46630;
	assign w11181 = w11106 ^ w11196;
	assign w11172 = w11196 & w11181;
	assign w11068 = w11108 ^ w11106;
	assign w11184 = w11105 ^ w11068;
	assign w11171 = w11193 & w11184;
	assign w11107 = w46634 ^ w11105;
	assign w11183 = w46630 ^ w11107;
	assign w11180 = w46631 ^ w11107;
	assign w11176 = w11195 & w11180;
	assign w11110 = w11176 ^ w11106;
	assign w11173 = w11194 & w11183;
	assign w11109 = w11173 ^ w11107;
	assign w11081 = w11172 ^ w11173;
	assign w11186 = w11105 ^ w11194;
	assign w11185 = w46636 ^ w11186;
	assign w11128 = w11081 ^ w11082;
	assign w11122 = w46635 ^ w46634;
	assign w11187 = w11122 ^ w11189;
	assign w11178 = w11187 & w11185;
	assign w11190 = w11194 ^ w11122;
	assign w11179 = w11186 & w11190;
	assign w11111 = w11179 ^ w11108;
	assign w11115 = w11111 ^ w11109;
	assign w11120 = w46629 ^ w11115;
	assign w11067 = w11108 ^ w46631;
	assign w11191 = w46636 ^ w11067;
	assign w11177 = w46636 & w11191;
	assign w43837 = w11171 ^ w11177;
	assign w11083 = w11115 ^ w43837;
	assign w11126 = w46631 ^ w11083;
	assign w11121 = w43837 ^ w11106;
	assign w11182 = w11112 ^ w11107;
	assign w11174 = w11189 & w11182;
	assign w43838 = w11171 ^ w11174;
	assign w11124 = w11172 ^ w43838;
	assign w11084 = w11110 ^ w43838;
	assign w11168 = w11084 ^ w11109;
	assign w11080 = w11175 ^ w11124;
	assign w11162 = w46635 ^ w11080;
	assign w11127 = w11128 ^ w11110;
	assign w11169 = w11175 ^ w11127;
	assign w11129 = w11172 ^ w11178;
	assign w11167 = w11129 ^ w11121;
	assign w11170 = w11129 ^ w11120;
	assign w11166 = w11170 & w11169;
	assign w11165 = w11166 ^ w11168;
	assign w11164 = w11167 & w11165;
	assign w11075 = w11164 ^ w11176;
	assign w11072 = w11164 ^ w11120;
	assign w11071 = w11075 ^ w11111;
	assign w11070 = w46631 ^ w11071;
	assign w11074 = w46629 ^ w11071;
	assign w11161 = w11166 ^ w11126;
	assign w11160 = w11161 & w11162;
	assign w11079 = w11160 ^ w11124;
	assign w11078 = w11160 ^ w11177;
	assign w11159 = w11160 ^ w11168;
	assign w11136 = w11159 & w11191;
	assign w11073 = w11078 ^ w11174;
	assign w11151 = w11073 ^ w11074;
	assign w11132 = w11151 & w11194;
	assign w11141 = w11151 & w11183;
	assign w11158 = w11166 ^ w11160;
	assign w11157 = w11168 & w11158;
	assign w43841 = w11157 ^ w11175;
	assign w11116 = w46635 ^ w43841;
	assign w11156 = w11116 ^ w11079;
	assign w11146 = w11156 & w11185;
	assign w11155 = w11157 ^ w11165;
	assign w11145 = w11159 & w46636;
	assign w11137 = w11156 & w11187;
	assign w11163 = w11164 ^ w11126;
	assign w11142 = w11163 & w11182;
	assign w11154 = w11163 & w11155;
	assign w11119 = w11154 ^ w11129;
	assign w11153 = w11119 ^ w11121;
	assign w11134 = w11153 & w11188;
	assign w11104 = w11142 ^ w11134;
	assign w11143 = w11153 & w11192;
	assign w11133 = w11163 & w11189;
	assign w11086 = w11142 ^ w11143;
	assign w11150 = w11119 ^ w11072;
	assign w11144 = w11150 & w11180;
	assign w43839 = w11143 ^ w11144;
	assign w11135 = w11150 & w11195;
	assign w11102 = w11144 ^ w11135;
	assign w11077 = w11154 ^ w11178;
	assign w11069 = w11116 ^ w11077;
	assign w11148 = w11069 ^ w11070;
	assign w11131 = w11148 & w11196;
	assign w43526 = w11131 ^ w11132;
	assign w11100 = w11104 ^ w43526;
	assign w11113 = w11137 ^ w43526;
	assign w11140 = w11148 & w11181;
	assign w11097 = w11140 ^ w11141;
	assign w11125 = w11140 ^ w43839;
	assign w11085 = w11141 ^ w11125;
	assign w11076 = w11106 ^ w11069;
	assign w11152 = w11073 ^ w11076;
	assign w11130 = w11152 & w11193;
	assign w11139 = w11152 & w11184;
	assign w11096 = w11141 ^ w11130;
	assign w11092 = ~w11096;
	assign w11091 = w11136 ^ w11125;
	assign w11088 = ~w11091;
	assign w11101 = w11140 ^ w11143;
	assign w11098 = ~w11101;
	assign w11117 = w11135 ^ w11139;
	assign w11095 = ~w11117;
	assign w11094 = w11095 ^ w11133;
	assign w11099 = w11095 ^ w11100;
	assign w11199 = w11098 ^ w11099;
	assign w50270 = ~w11199;
	assign w43460 = w45586 ^ w50270;
	assign w43176 = w11199 ^ w45587;
	assign w43509 = w43175 ^ w43176;
	assign w11149 = w43841 ^ w11127;
	assign w11138 = w11149 & w11190;
	assign w11147 = w11149 & w11186;
	assign w11114 = w11138 ^ w11113;
	assign w50274 = w11114 ^ w11085;
	assign w43421 = w50269 ^ w50274;
	assign w43284 = w43421 ^ w45674;
	assign w43840 = w11145 ^ w11147;
	assign w11103 = w43840 ^ w11100;
	assign w11200 = w11102 ^ w11103;
	assign w11090 = w11094 ^ w43840;
	assign w11089 = w11113 ^ w11090;
	assign w50271 = w11088 ^ w11089;
	assign w43456 = w50266 ^ w50271;
	assign w43335 = w50271 ^ w45586;
	assign w43309 = ~w43456;
	assign w43307 = w43309 ^ w50279;
	assign w11118 = w11146 ^ w11114;
	assign w11123 = w11147 ^ w11118;
	assign w11198 = w11123 ^ w11097;
	assign w11087 = w11145 ^ w11118;
	assign w50272 = w11086 ^ w11087;
	assign w43453 = w50267 ^ w50272;
	assign w43317 = ~w43453;
	assign w43180 = ~w50272;
	assign w43179 = w43180 ^ w50266;
	assign w43508 = w43178 ^ w43179;
	assign w45222 = ~w11198;
	assign w45223 = ~w11200;
	assign w43461 = w45587 ^ w45223;
	assign w50273 = w43839 ^ w11123;
	assign w43449 = w50268 ^ w50273;
	assign w43291 = ~w43449;
	assign w43182 = w50273 ^ w50267;
	assign w43507 = w43181 ^ w43182;
	assign w11093 = w11132 ^ w11090;
	assign w11197 = w11092 ^ w11093;
	assign w45229 = ~w11197;
	assign w43445 = w45592 ^ w45229;
	assign w43333 = w45229 ^ w50268;
	assign w43313 = w43445 ^ w43439;
	assign w43306 = w43445 ^ w45681;
	assign w43304 = ~w43306;
	assign w43303 = w45222 ^ w45229;
	assign w45949 = ~w9485;
	assign w9430 = w45949 ^ w50047;
	assign w49929 = w9429 ^ w9430;
	assign w9409 = w45949 ^ w50064;
	assign w49940 = w9409 ^ w9410;
	assign w46728 = w49929 ^ w1194;
	assign w46717 = w49940 ^ w1205;
	assign w26650 = w46719 ^ w46717;
	assign w26612 = w26652 ^ w26650;
	assign w26728 = w26649 ^ w26612;
	assign w9273 = w45949 ^ w45766;
	assign w11376 = w46728 ^ w46726;
	assign w11335 = w11376 ^ w46727;
	assign w11336 = w11376 ^ w11374;
	assign w26725 = w26650 ^ w26740;
	assign w11462 = w46728 ^ w46725;
	assign w26716 = w26740 & w26725;
	assign w26739 = w46717 ^ w46723;
	assign w26720 = w26739 & w26724;
	assign w26654 = w26720 ^ w26650;
	assign w9555 = w9273 ^ w9274;
	assign w49926 = w9555 ^ w9547;
	assign w46731 = w49926 ^ w1191;
	assign w11456 = w46731 ^ w11460;
	assign w11390 = w46731 ^ w46730;
	assign w11455 = w11390 ^ w11457;
	assign w11443 = w11460 & w11456;
	assign w11373 = w46731 ^ w46729;
	assign w11454 = w11373 ^ w11462;
	assign w11375 = w46730 ^ w11373;
	assign w11448 = w46727 ^ w11375;
	assign w11450 = w11380 ^ w11375;
	assign w11451 = w46726 ^ w11375;
	assign w11453 = w46732 ^ w11454;
	assign w11441 = w11462 & w11451;
	assign w11377 = w11441 ^ w11375;
	assign w11463 = w46725 ^ w46731;
	assign w11444 = w11463 & w11448;
	assign w11378 = w11444 ^ w11374;
	assign w11452 = w11373 ^ w11336;
	assign w11439 = w11461 & w11452;
	assign w11442 = w11457 & w11450;
	assign w43849 = w11439 ^ w11442;
	assign w11352 = w11378 ^ w43849;
	assign w11436 = w11352 ^ w11377;
	assign w11459 = w46732 ^ w11335;
	assign w11445 = w46732 & w11459;
	assign w43848 = w11439 ^ w11445;
	assign w11389 = w43848 ^ w11374;
	assign w26738 = w46720 ^ w46717;
	assign w26730 = w26649 ^ w26738;
	assign w26734 = w26738 ^ w26666;
	assign w26723 = w26730 & w26734;
	assign w26655 = w26723 ^ w26652;
	assign w26717 = w26738 & w26727;
	assign w26653 = w26717 ^ w26651;
	assign w26659 = w26655 ^ w26653;
	assign w26625 = w26716 ^ w26717;
	assign w26672 = w26625 ^ w26626;
	assign w26671 = w26672 ^ w26654;
	assign w26713 = w26719 ^ w26671;
	assign w26737 = w46717 ^ w46722;
	assign w26715 = w26737 & w26728;
	assign w44485 = w26715 ^ w26721;
	assign w26665 = w44485 ^ w26650;
	assign w11464 = w46730 ^ w46728;
	assign w11449 = w11374 ^ w11464;
	assign w11440 = w11464 & w11449;
	assign w11349 = w11440 ^ w11441;
	assign w11396 = w11349 ^ w11350;
	assign w11395 = w11396 ^ w11378;
	assign w11437 = w11443 ^ w11395;
	assign w11392 = w11440 ^ w43849;
	assign w11348 = w11443 ^ w11392;
	assign w11430 = w46731 ^ w11348;
	assign w11446 = w11455 & w11453;
	assign w11397 = w11440 ^ w11446;
	assign w11435 = w11397 ^ w11389;
	assign w26733 = w26650 ^ w26656;
	assign w26718 = w26733 & w26726;
	assign w26731 = w26666 ^ w26733;
	assign w44486 = w26715 ^ w26718;
	assign w26628 = w26654 ^ w44486;
	assign w26712 = w26628 ^ w26653;
	assign w26668 = w26716 ^ w44486;
	assign w26624 = w26719 ^ w26668;
	assign w26706 = w46723 ^ w26624;
	assign w11458 = w11462 ^ w11390;
	assign w11447 = w11454 & w11458;
	assign w11379 = w11447 ^ w11376;
	assign w11383 = w11379 ^ w11377;
	assign w11351 = w11383 ^ w43848;
	assign w11394 = w46727 ^ w11351;
	assign w11388 = w46725 ^ w11383;
	assign w11438 = w11397 ^ w11388;
	assign w11434 = w11438 & w11437;
	assign w11429 = w11434 ^ w11394;
	assign w11428 = w11429 & w11430;
	assign w11426 = w11434 ^ w11428;
	assign w11427 = w11428 ^ w11436;
	assign w11404 = w11427 & w11459;
	assign w11413 = w11427 & w46732;
	assign w11347 = w11428 ^ w11392;
	assign w11346 = w11428 ^ w11445;
	assign w11425 = w11436 & w11426;
	assign w11341 = w11346 ^ w11442;
	assign w43852 = w11425 ^ w11443;
	assign w11384 = w46731 ^ w43852;
	assign w11424 = w11384 ^ w11347;
	assign w11414 = w11424 & w11453;
	assign w11405 = w11424 & w11455;
	assign w11417 = w43852 ^ w11395;
	assign w11415 = w11417 & w11454;
	assign w11406 = w11417 & w11458;
	assign w43851 = w11413 ^ w11415;
	assign w11433 = w11434 ^ w11436;
	assign w11423 = w11425 ^ w11433;
	assign w11432 = w11435 & w11433;
	assign w11431 = w11432 ^ w11394;
	assign w11401 = w11431 & w11457;
	assign w11422 = w11431 & w11423;
	assign w11387 = w11422 ^ w11397;
	assign w11345 = w11422 ^ w11446;
	assign w11337 = w11384 ^ w11345;
	assign w11421 = w11387 ^ w11389;
	assign w11402 = w11421 & w11456;
	assign w11344 = w11374 ^ w11337;
	assign w11340 = w11432 ^ w11388;
	assign w11418 = w11387 ^ w11340;
	assign w11403 = w11418 & w11463;
	assign w11343 = w11432 ^ w11444;
	assign w11412 = w11418 & w11448;
	assign w11370 = w11412 ^ w11403;
	assign w11339 = w11343 ^ w11379;
	assign w11342 = w46725 ^ w11339;
	assign w11419 = w11341 ^ w11342;
	assign w11400 = w11419 & w11462;
	assign w11409 = w11419 & w11451;
	assign w11410 = w11431 & w11450;
	assign w11372 = w11410 ^ w11402;
	assign w11411 = w11421 & w11460;
	assign w11354 = w11410 ^ w11411;
	assign w43850 = w11411 ^ w11412;
	assign w11420 = w11341 ^ w11344;
	assign w11407 = w11420 & w11452;
	assign w11398 = w11420 & w11461;
	assign w11385 = w11403 ^ w11407;
	assign w11364 = w11409 ^ w11398;
	assign w11360 = ~w11364;
	assign w11338 = w46727 ^ w11339;
	assign w11416 = w11337 ^ w11338;
	assign w11399 = w11416 & w11464;
	assign w43527 = w11399 ^ w11400;
	assign w11368 = w11372 ^ w43527;
	assign w11371 = w43851 ^ w11368;
	assign w11468 = w11370 ^ w11371;
	assign w11381 = w11405 ^ w43527;
	assign w11382 = w11406 ^ w11381;
	assign w11386 = w11414 ^ w11382;
	assign w11355 = w11413 ^ w11386;
	assign w50289 = w11354 ^ w11355;
	assign w11391 = w11415 ^ w11386;
	assign w50290 = w43850 ^ w11391;
	assign w43462 = w50285 ^ w50290;
	assign w43470 = w50284 ^ w50289;
	assign w43237 = ~w43470;
	assign w43260 = w43237 ^ w43450;
	assign w43259 = w43462 ^ w43444;
	assign w50195 = w45312 ^ w43259;
	assign w46535 = w50195 ^ w1258;
	assign w43250 = w50296 ^ w50290;
	assign w43235 = w43237 ^ w43469;
	assign w43234 = ~w43462;
	assign w43232 = w43234 ^ w43459;
	assign w43199 = ~w50289;
	assign w43209 = w50295 ^ w43199;
	assign w43201 = w50290 ^ w50284;
	assign w43499 = w43200 ^ w43201;
	assign w50186 = w43499 ^ w43450;
	assign w46544 = w50186 ^ w1249;
	assign w43198 = w43199 ^ w50283;
	assign w43500 = w43197 ^ w43198;
	assign w50185 = w43500 ^ w43459;
	assign w46545 = w50185 ^ w1248;
	assign w11408 = w11416 & w11449;
	assign w11393 = w11408 ^ w43850;
	assign w11353 = w11409 ^ w11393;
	assign w50293 = w11382 ^ w11353;
	assign w43422 = w50286 ^ w50293;
	assign w43426 = w50293 ^ w50297;
	assign w43270 = w50293 ^ w45313;
	assign w50189 = w43269 ^ w43270;
	assign w46541 = w50189 ^ w1252;
	assign w43268 = w43481 ^ w43422;
	assign w50190 = w45307 ^ w43268;
	assign w46540 = w50190 ^ w1253;
	assign w43229 = w43433 ^ w43422;
	assign w50213 = w50297 ^ w43229;
	assign w43207 = ~w43426;
	assign w43208 = w43207 ^ w50300;
	assign w43496 = w43208 ^ w43209;
	assign w50202 = w43496 ^ w43462;
	assign w46528 = w50202 ^ w1265;
	assign w43204 = w43207 ^ w50299;
	assign w43202 = w43426 ^ w45511;
	assign w46517 = w50213 ^ w1276;
	assign w45226 = ~w11468;
	assign w43485 = w45307 ^ w45226;
	assign w50182 = w45226 ^ w43283;
	assign w46548 = w50182 ^ w1245;
	assign w43266 = w43485 ^ w43473;
	assign w43254 = w43485 ^ w43426;
	assign w50198 = w45512 ^ w43254;
	assign w46532 = w50198 ^ w1261;
	assign w43243 = w43485 ^ w43419;
	assign w50206 = w45315 ^ w43243;
	assign w46524 = w50206 ^ w1269;
	assign w43203 = w45315 ^ w45226;
	assign w43498 = w43202 ^ w43203;
	assign w11359 = w11404 ^ w11393;
	assign w11356 = ~w11359;
	assign w11369 = w11408 ^ w11411;
	assign w11366 = ~w11369;
	assign w45898 = ~w43422;
	assign w43267 = w45898 ^ w45306;
	assign w43265 = w43266 ^ w43267;
	assign w50191 = ~w43265;
	assign w43263 = w45898 ^ w50284;
	assign w43261 = w45898 ^ w50285;
	assign w50194 = w43260 ^ w43261;
	assign w46536 = w50194 ^ w1257;
	assign w43244 = w45898 ^ w50301;
	assign w46539 = w50191 ^ w1254;
	assign w26729 = w46724 ^ w26730;
	assign w26722 = w26731 & w26729;
	assign w26673 = w26716 ^ w26722;
	assign w26711 = w26673 ^ w26665;
	assign w11363 = ~w11385;
	assign w11367 = w11363 ^ w11368;
	assign w11467 = w11366 ^ w11367;
	assign w50287 = ~w11467;
	assign w43484 = w45306 ^ w50287;
	assign w50199 = w43498 ^ w43484;
	assign w46531 = w50199 ^ w1262;
	assign w43264 = w43484 ^ w43469;
	assign w50192 = w50283 ^ w43264;
	assign w46538 = w50192 ^ w1255;
	assign w10854 = w46539 ^ w46538;
	assign w43252 = w45314 ^ w11467;
	assign w43242 = w43484 ^ w43481;
	assign w43240 = ~w43242;
	assign w43195 = w11467 ^ w45307;
	assign w43501 = w43194 ^ w43195;
	assign w50183 = w43501 ^ w43473;
	assign w46547 = w50183 ^ w1246;
	assign w14589 = w46547 ^ w46545;
	assign w14679 = w46541 ^ w46547;
	assign w10928 = w46538 ^ w46536;
	assign w11362 = w11363 ^ w11401;
	assign w11358 = w11362 ^ w43851;
	assign w11361 = w11400 ^ w11358;
	assign w11465 = w11360 ^ w11361;
	assign w50291 = ~w11465;
	assign w43455 = w45312 ^ w50291;
	assign w43278 = w11465 ^ w50285;
	assign w50187 = w43277 ^ w43278;
	assign w46543 = w50187 ^ w1250;
	assign w14590 = w46543 ^ w46541;
	assign w43258 = w43455 ^ w43433;
	assign w50196 = w45313 ^ w43258;
	assign w46534 = w50196 ^ w1259;
	assign w43249 = w43455 ^ w45517;
	assign w50203 = w43249 ^ w43250;
	assign w46527 = w50203 ^ w1266;
	assign w43247 = w45320 ^ w11465;
	assign w43231 = w43455 ^ w43450;
	assign w50211 = w45320 ^ w43231;
	assign w46519 = w50211 ^ w1274;
	assign w10840 = w46536 ^ w46534;
	assign w10799 = w10840 ^ w46535;
	assign w10923 = w46540 ^ w10799;
	assign w29196 = w46519 ^ w46517;
	assign w10909 = w46540 & w10923;
	assign w11357 = w11381 ^ w11358;
	assign w50288 = w11356 ^ w11357;
	assign w43477 = w50283 ^ w50288;
	assign w43206 = ~w50288;
	assign w43281 = w43206 ^ w45306;
	assign w50184 = w43280 ^ w43281;
	assign w46546 = w50184 ^ w1247;
	assign w14606 = w46547 ^ w46546;
	assign w14680 = w46546 ^ w46544;
	assign w14591 = w46546 ^ w14589;
	assign w14664 = w46543 ^ w14591;
	assign w14660 = w14679 & w14664;
	assign w14594 = w14660 ^ w14590;
	assign w14665 = w14590 ^ w14680;
	assign w14656 = w14680 & w14665;
	assign w43253 = ~w43477;
	assign w43262 = w43253 ^ w43459;
	assign w50193 = w43262 ^ w43263;
	assign w46537 = w50193 ^ w1256;
	assign w10837 = w46539 ^ w46537;
	assign w43251 = w43253 ^ w50298;
	assign w50200 = w43251 ^ w43252;
	assign w46530 = w50200 ^ w1263;
	assign w26204 = w46530 ^ w46528;
	assign w43238 = w43477 ^ w43473;
	assign w50208 = w50294 ^ w43238;
	assign w43205 = w50294 ^ w43206;
	assign w43497 = w43204 ^ w43205;
	assign w50201 = w43497 ^ w43470;
	assign w10814 = w46537 ^ w46538;
	assign w46522 = w50208 ^ w1271;
	assign w29283 = w46517 ^ w46522;
	assign w10839 = w46538 ^ w10837;
	assign w10915 = w46534 ^ w10839;
	assign w10912 = w46535 ^ w10839;
	assign w26130 = w46531 ^ w46530;
	assign w14677 = w46541 ^ w46546;
	assign w14566 = w46545 ^ w46546;
	assign w46529 = w50201 ^ w1264;
	assign w26113 = w46531 ^ w46529;
	assign w26115 = w46530 ^ w26113;
	assign w26188 = w46527 ^ w26115;
	assign w26090 = w46529 ^ w46530;
	assign w26627 = w26659 ^ w44485;
	assign w26670 = w46719 ^ w26627;
	assign w26664 = w46717 ^ w26659;
	assign w26714 = w26673 ^ w26664;
	assign w26710 = w26714 & w26713;
	assign w26709 = w26710 ^ w26712;
	assign w26708 = w26711 & w26709;
	assign w26616 = w26708 ^ w26664;
	assign w26707 = w26708 ^ w26670;
	assign w26677 = w26707 & w26733;
	assign w26705 = w26710 ^ w26670;
	assign w26704 = w26705 & w26706;
	assign w26623 = w26704 ^ w26668;
	assign w26702 = w26710 ^ w26704;
	assign w26703 = w26704 ^ w26712;
	assign w26701 = w26712 & w26702;
	assign w26699 = w26701 ^ w26709;
	assign w26698 = w26707 & w26699;
	assign w26680 = w26703 & w26735;
	assign w26686 = w26707 & w26726;
	assign w44489 = w26701 ^ w26719;
	assign w26693 = w44489 ^ w26671;
	assign w26682 = w26693 & w26734;
	assign w26691 = w26693 & w26730;
	assign w26621 = w26698 ^ w26722;
	assign w26660 = w46723 ^ w44489;
	assign w26700 = w26660 ^ w26623;
	assign w26690 = w26700 & w26729;
	assign w26681 = w26700 & w26731;
	assign w26613 = w26660 ^ w26621;
	assign w26620 = w26650 ^ w26613;
	assign w26619 = w26708 ^ w26720;
	assign w26615 = w26619 ^ w26655;
	assign w26614 = w46719 ^ w26615;
	assign w26692 = w26613 ^ w26614;
	assign w26684 = w26692 & w26725;
	assign w26618 = w46717 ^ w26615;
	assign w26675 = w26692 & w26740;
	assign w26689 = w26703 & w46724;
	assign w44488 = w26689 ^ w26691;
	assign w26663 = w26698 ^ w26673;
	assign w26694 = w26663 ^ w26616;
	assign w26697 = w26663 ^ w26665;
	assign w26687 = w26697 & w26736;
	assign w26645 = w26684 ^ w26687;
	assign w26642 = ~w26645;
	assign w26630 = w26686 ^ w26687;
	assign w26679 = w26694 & w26739;
	assign w26622 = w26704 ^ w26721;
	assign w26617 = w26622 ^ w26718;
	assign w26695 = w26617 ^ w26618;
	assign w26696 = w26617 ^ w26620;
	assign w26683 = w26696 & w26728;
	assign w26661 = w26679 ^ w26683;
	assign w26674 = w26696 & w26737;
	assign w26639 = ~w26661;
	assign w26638 = w26639 ^ w26677;
	assign w26685 = w26695 & w26727;
	assign w26640 = w26685 ^ w26674;
	assign w26634 = w26638 ^ w44488;
	assign w26641 = w26684 ^ w26685;
	assign w26676 = w26695 & w26738;
	assign w26637 = w26676 ^ w26634;
	assign w43574 = w26675 ^ w26676;
	assign w26657 = w26681 ^ w43574;
	assign w26633 = w26657 ^ w26634;
	assign w26658 = w26682 ^ w26657;
	assign w26662 = w26690 ^ w26658;
	assign w26631 = w26689 ^ w26662;
	assign w50276 = w26630 ^ w26631;
	assign w43446 = w50276 ^ w50280;
	assign w50153 = w43508 ^ w43446;
	assign w46577 = w50153 ^ w1280;
	assign w43318 = w43309 ^ w43446;
	assign w43288 = w43291 ^ w43446;
	assign w43192 = w50276 ^ w43180;
	assign w26667 = w26691 ^ w26662;
	assign w26742 = w26667 ^ w26641;
	assign w26636 = ~w26640;
	assign w26741 = w26636 ^ w26637;
	assign w26688 = w26694 & w26724;
	assign w26646 = w26688 ^ w26679;
	assign w44487 = w26687 ^ w26688;
	assign w50277 = w44487 ^ w26667;
	assign w43441 = w50277 ^ w50281;
	assign w50154 = w43507 ^ w43441;
	assign w46576 = w50154 ^ w1281;
	assign w43315 = w43317 ^ w43441;
	assign w43290 = ~w50277;
	assign w43305 = w43290 ^ w50273;
	assign w50171 = w43304 ^ w43305;
	assign w43287 = w43445 ^ w43441;
	assign w26669 = w26684 ^ w44487;
	assign w26629 = w26685 ^ w26669;
	assign w50278 = w26658 ^ w26629;
	assign w43420 = w50278 ^ w50282;
	assign w43428 = w50274 ^ w50278;
	assign w43329 = w43439 ^ w43420;
	assign w50157 = w50274 ^ w43329;
	assign w46573 = w50157 ^ w1284;
	assign w26336 = w46576 ^ w46573;
	assign w43311 = w43420 ^ w45222;
	assign w50165 = w43311 ^ w43312;
	assign w46565 = w50165 ^ w1292;
	assign w43310 = w43461 ^ w43428;
	assign w50166 = w45676 ^ w43310;
	assign w46564 = w50166 ^ w1293;
	assign w43300 = w43461 ^ w43420;
	assign w43296 = w43420 ^ w50276;
	assign w43289 = w43420 ^ w43290;
	assign w50178 = w43288 ^ w43289;
	assign w46552 = w50178 ^ w1305;
	assign w43193 = ~w43428;
	assign w43191 = w43193 ^ w50281;
	assign w43502 = w43191 ^ w43192;
	assign w50170 = w43502 ^ w43449;
	assign w46560 = w50170 ^ w1297;
	assign w43189 = w43428 ^ w50280;
	assign w43187 = w43428 ^ w45675;
	assign w26635 = w26680 ^ w26669;
	assign w26632 = ~w26635;
	assign w50275 = w26632 ^ w26633;
	assign w43451 = w50275 ^ w50279;
	assign w43334 = w43451 ^ w45675;
	assign w50152 = w43334 ^ w43335;
	assign w46578 = w50152 ^ w1279;
	assign w26224 = w46577 ^ w46578;
	assign w26338 = w46578 ^ w46576;
	assign w43320 = w43460 ^ w43451;
	assign w50160 = w50266 ^ w43320;
	assign w46570 = w50160 ^ w1287;
	assign w11059 = w46565 ^ w46570;
	assign w43295 = w43453 ^ w43451;
	assign w50177 = w43295 ^ w43296;
	assign w46553 = w50177 ^ w1304;
	assign w43190 = w50275 ^ w50271;
	assign w43503 = w43189 ^ w43190;
	assign w50169 = w43503 ^ w43453;
	assign w46559 = w50171 ^ w1298;
	assign w46561 = w50169 ^ w1296;
	assign w26335 = w46573 ^ w46578;
	assign w45596 = ~w26741;
	assign w43436 = w45596 ^ w45681;
	assign w43332 = w43436 ^ w50281;
	assign w50155 = w43332 ^ w43333;
	assign w43314 = w43449 ^ w43436;
	assign w50163 = w45592 ^ w43314;
	assign w46567 = w50163 ^ w1290;
	assign w10972 = w46567 ^ w46565;
	assign w43302 = w43439 ^ w45596;
	assign w50172 = w43302 ^ w43303;
	assign w46558 = w50172 ^ w1299;
	assign w14730 = w46564 ^ w46558;
	assign w14810 = w46559 ^ w14730;
	assign w50179 = w45596 ^ w43287;
	assign w46551 = w50179 ^ w1306;
	assign w46575 = w50155 ^ w1282;
	assign w26248 = w46575 ^ w46573;
	assign w26323 = w26248 ^ w26338;
	assign w14726 = w46560 ^ w46558;
	assign w14685 = w14726 ^ w46559;
	assign w26314 = w26338 & w26323;
	assign w14809 = w46564 ^ w14685;
	assign w14795 = w46564 & w14809;
	assign w45597 = ~w26742;
	assign w43438 = w45222 ^ w45597;
	assign w43330 = w43438 ^ w45674;
	assign w50156 = w43330 ^ w43331;
	assign w46574 = w50156 ^ w1283;
	assign w50164 = w45597 ^ w43313;
	assign w46566 = w50164 ^ w1291;
	assign w43301 = w43438 ^ w43421;
	assign w50173 = w50282 ^ w43301;
	assign w43286 = w43438 ^ w43436;
	assign w50180 = w45593 ^ w43286;
	assign w46550 = w50180 ^ w1307;
	assign w23570 = w46552 ^ w46550;
	assign w43285 = w50278 ^ w45597;
	assign w50181 = w43284 ^ w43285;
	assign w46549 = w50181 ^ w1308;
	assign w23656 = w46552 ^ w46549;
	assign w23568 = w46551 ^ w46549;
	assign w23530 = w23570 ^ w23568;
	assign w23529 = w23570 ^ w46551;
	assign w26250 = w46576 ^ w46574;
	assign w26210 = w26250 ^ w26248;
	assign w26209 = w26250 ^ w46575;
	assign w46557 = w50173 ^ w1300;
	assign w14724 = w46559 ^ w46557;
	assign w14807 = w14724 ^ w14730;
	assign w14812 = w46560 ^ w46557;
	assign w14686 = w14726 ^ w14724;
	assign w26678 = w26697 & w26732;
	assign w26648 = w26686 ^ w26678;
	assign w26644 = w26648 ^ w43574;
	assign w26643 = w26639 ^ w26644;
	assign w26743 = w26642 ^ w26643;
	assign w26647 = w44488 ^ w26644;
	assign w26744 = w26646 ^ w26647;
	assign w45590 = ~w26743;
	assign w43454 = w45590 ^ w45675;
	assign w50151 = w43509 ^ w43454;
	assign w46579 = w50151 ^ w1278;
	assign w26337 = w46573 ^ w46579;
	assign w26247 = w46579 ^ w46577;
	assign w26249 = w46578 ^ w26247;
	assign w26322 = w46575 ^ w26249;
	assign w26318 = w26337 & w26322;
	assign w26325 = w46574 ^ w26249;
	assign w43322 = w43461 ^ w43454;
	assign w43308 = w45590 ^ w11199;
	assign w50168 = w43307 ^ w43308;
	assign w46562 = w50168 ^ w1295;
	assign w14811 = w46557 ^ w46562;
	assign w14814 = w46562 ^ w46560;
	assign w14799 = w14724 ^ w14814;
	assign w14700 = w46561 ^ w46562;
	assign w43299 = w43420 ^ w45590;
	assign w43297 = w43456 ^ w43454;
	assign w50176 = w50275 ^ w43297;
	assign w46554 = w50176 ^ w1303;
	assign w23544 = w46553 ^ w46554;
	assign w26264 = w46579 ^ w46578;
	assign w26332 = w26336 ^ w26264;
	assign w26326 = w26247 ^ w26210;
	assign w26313 = w26335 & w26326;
	assign w23658 = w46554 ^ w46552;
	assign w26252 = w26318 ^ w26248;
	assign w26315 = w26336 & w26325;
	assign w26223 = w26314 ^ w26315;
	assign w26251 = w26315 ^ w26249;
	assign w23655 = w46549 ^ w46554;
	assign w26328 = w26247 ^ w26336;
	assign w26321 = w26328 & w26332;
	assign w26253 = w26321 ^ w26250;
	assign w26257 = w26253 ^ w26251;
	assign w26262 = w46573 ^ w26257;
	assign w14790 = w14814 & w14799;
	assign w45591 = ~w26744;
	assign w43458 = w45591 ^ w45676;
	assign w43336 = w43458 ^ w43430;
	assign w50150 = w45223 ^ w43336;
	assign w46580 = w50150 ^ w1277;
	assign w26333 = w46580 ^ w26209;
	assign w26327 = w46580 ^ w26328;
	assign w43324 = w43458 ^ w43421;
	assign w50158 = w45587 ^ w43324;
	assign w46572 = w50158 ^ w1285;
	assign w10978 = w46572 ^ w46566;
	assign w11055 = w10972 ^ w10978;
	assign w50174 = w45591 ^ w43300;
	assign w46556 = w50174 ^ w1301;
	assign w43298 = w43460 ^ w43458;
	assign w50175 = w43298 ^ w43299;
	assign w46555 = w50175 ^ w1302;
	assign w23657 = w46549 ^ w46555;
	assign w23567 = w46555 ^ w46553;
	assign w23648 = w23567 ^ w23656;
	assign w23646 = w23567 ^ w23530;
	assign w23633 = w23655 & w23646;
	assign w23569 = w46554 ^ w23567;
	assign w43188 = w45591 ^ w45223;
	assign w43504 = w43187 ^ w43188;
	assign w50167 = w43504 ^ w43460;
	assign w46563 = w50167 ^ w1294;
	assign w14806 = w46563 ^ w14810;
	assign w14740 = w46563 ^ w46562;
	assign w14805 = w14740 ^ w14807;
	assign w14808 = w14812 ^ w14740;
	assign w14813 = w46557 ^ w46563;
	assign w23653 = w46556 ^ w23529;
	assign w14723 = w46563 ^ w46561;
	assign w14804 = w14723 ^ w14812;
	assign w14803 = w46564 ^ w14804;
	assign w14796 = w14805 & w14803;
	assign w14797 = w14804 & w14808;
	assign w26319 = w46580 & w26333;
	assign w44471 = w26313 ^ w26319;
	assign w26225 = w26257 ^ w44471;
	assign w26268 = w46575 ^ w26225;
	assign w23645 = w46550 ^ w23569;
	assign w23574 = w46556 ^ w46550;
	assign w23651 = w23568 ^ w23574;
	assign w23644 = w23574 ^ w23569;
	assign w23647 = w46556 ^ w23648;
	assign w26254 = w46580 ^ w46574;
	assign w26324 = w26254 ^ w26249;
	assign w23636 = w23651 & w23644;
	assign w44357 = w23633 ^ w23636;
	assign w26331 = w26248 ^ w26254;
	assign w26329 = w26264 ^ w26331;
	assign w26320 = w26329 & w26327;
	assign w26316 = w26331 & w26324;
	assign w44468 = w26313 ^ w26316;
	assign w26226 = w26252 ^ w44468;
	assign w26310 = w26226 ^ w26251;
	assign w14747 = w14790 ^ w14796;
	assign w11058 = w46567 ^ w10978;
	assign w14793 = w14810 & w14806;
	assign w23654 = w46551 ^ w23574;
	assign w23650 = w46555 ^ w23654;
	assign w14725 = w46562 ^ w14723;
	assign w14798 = w46559 ^ w14725;
	assign w14794 = w14813 & w14798;
	assign w14728 = w14794 ^ w14724;
	assign w14801 = w46558 ^ w14725;
	assign w14800 = w14730 ^ w14725;
	assign w14792 = w14807 & w14800;
	assign w26263 = w44471 ^ w26248;
	assign w26266 = w26314 ^ w44468;
	assign w26271 = w26314 ^ w26320;
	assign w26309 = w26271 ^ w26263;
	assign w26312 = w26271 ^ w26262;
	assign w14729 = w14797 ^ w14726;
	assign w23639 = w46556 & w23653;
	assign w44360 = w23633 ^ w23639;
	assign w23583 = w44360 ^ w23568;
	assign w23637 = w23654 & w23650;
	assign w23635 = w23656 & w23645;
	assign w23571 = w23635 ^ w23569;
	assign w14791 = w14812 & w14801;
	assign w14727 = w14791 ^ w14725;
	assign w14699 = w14790 ^ w14791;
	assign w14746 = w14699 ^ w14700;
	assign w14745 = w14746 ^ w14728;
	assign w14733 = w14729 ^ w14727;
	assign w14738 = w46557 ^ w14733;
	assign w14788 = w14747 ^ w14738;
	assign w14787 = w14793 ^ w14745;
	assign w14784 = w14788 & w14787;
	assign w23642 = w46551 ^ w23569;
	assign w23638 = w23657 & w23642;
	assign w23572 = w23638 ^ w23568;
	assign w23643 = w23568 ^ w23658;
	assign w23634 = w23658 & w23643;
	assign w23543 = w23634 ^ w23635;
	assign w23590 = w23543 ^ w23544;
	assign w23586 = w23634 ^ w44357;
	assign w23542 = w23637 ^ w23586;
	assign w23624 = w46555 ^ w23542;
	assign w23589 = w23590 ^ w23572;
	assign w23631 = w23637 ^ w23589;
	assign w14802 = w14723 ^ w14686;
	assign w14789 = w14811 & w14802;
	assign w43987 = w14789 ^ w14795;
	assign w14739 = w43987 ^ w14724;
	assign w14785 = w14747 ^ w14739;
	assign w14701 = w14733 ^ w43987;
	assign w14744 = w46559 ^ w14701;
	assign w14779 = w14784 ^ w14744;
	assign w43988 = w14789 ^ w14792;
	assign w14742 = w14790 ^ w43988;
	assign w14698 = w14793 ^ w14742;
	assign w14780 = w46563 ^ w14698;
	assign w14702 = w14728 ^ w43988;
	assign w14786 = w14702 ^ w14727;
	assign w14778 = w14779 & w14780;
	assign w14776 = w14784 ^ w14778;
	assign w14696 = w14778 ^ w14795;
	assign w14777 = w14778 ^ w14786;
	assign w14763 = w14777 & w46564;
	assign w14697 = w14778 ^ w14742;
	assign w14775 = w14786 & w14776;
	assign w43991 = w14775 ^ w14793;
	assign w14767 = w43991 ^ w14745;
	assign w14765 = w14767 & w14804;
	assign w14756 = w14767 & w14808;
	assign w43990 = w14763 ^ w14765;
	assign w14734 = w46563 ^ w43991;
	assign w14774 = w14734 ^ w14697;
	assign w14764 = w14774 & w14803;
	assign w14755 = w14774 & w14805;
	assign w14754 = w14777 & w14809;
	assign w14783 = w14784 ^ w14786;
	assign w14782 = w14785 & w14783;
	assign w14693 = w14782 ^ w14794;
	assign w14689 = w14693 ^ w14729;
	assign w14692 = w46557 ^ w14689;
	assign w14690 = w14782 ^ w14738;
	assign w14781 = w14782 ^ w14744;
	assign w14751 = w14781 & w14807;
	assign w14773 = w14775 ^ w14783;
	assign w14760 = w14781 & w14800;
	assign w14688 = w46559 ^ w14689;
	assign w14691 = w14696 ^ w14792;
	assign w14769 = w14691 ^ w14692;
	assign w14750 = w14769 & w14812;
	assign w14759 = w14769 & w14801;
	assign w14772 = w14781 & w14773;
	assign w14737 = w14772 ^ w14747;
	assign w14771 = w14737 ^ w14739;
	assign w14752 = w14771 & w14806;
	assign w14722 = w14760 ^ w14752;
	assign w14761 = w14771 & w14810;
	assign w14768 = w14737 ^ w14690;
	assign w14753 = w14768 & w14813;
	assign w14762 = w14768 & w14798;
	assign w14720 = w14762 ^ w14753;
	assign w14695 = w14772 ^ w14796;
	assign w14687 = w14734 ^ w14695;
	assign w14694 = w14724 ^ w14687;
	assign w14770 = w14691 ^ w14694;
	assign w14757 = w14770 & w14802;
	assign w14735 = w14753 ^ w14757;
	assign w14713 = ~w14735;
	assign w14712 = w14713 ^ w14751;
	assign w14708 = w14712 ^ w43990;
	assign w43989 = w14761 ^ w14762;
	assign w14711 = w14750 ^ w14708;
	assign w14748 = w14770 & w14811;
	assign w14714 = w14759 ^ w14748;
	assign w14710 = ~w14714;
	assign w14815 = w14710 ^ w14711;
	assign w14766 = w14687 ^ w14688;
	assign w14749 = w14766 & w14814;
	assign w43538 = w14749 ^ w14750;
	assign w14731 = w14755 ^ w43538;
	assign w14707 = w14731 ^ w14708;
	assign w14718 = w14722 ^ w43538;
	assign w14721 = w43990 ^ w14718;
	assign w14818 = w14720 ^ w14721;
	assign w14717 = w14713 ^ w14718;
	assign w14758 = w14766 & w14799;
	assign w14715 = w14758 ^ w14759;
	assign w14719 = w14758 ^ w14761;
	assign w14716 = ~w14719;
	assign w14817 = w14716 ^ w14717;
	assign w14743 = w14758 ^ w43989;
	assign w14703 = w14759 ^ w14743;
	assign w14709 = w14754 ^ w14743;
	assign w14706 = ~w14709;
	assign w50495 = w14706 ^ w14707;
	assign w45294 = ~w14818;
	assign w45299 = ~w14815;
	assign w45301 = ~w14817;
	assign w14732 = w14756 ^ w14731;
	assign w50498 = w14732 ^ w14703;
	assign w14736 = w14764 ^ w14732;
	assign w14741 = w14765 ^ w14736;
	assign w50497 = w43989 ^ w14741;
	assign w14705 = w14763 ^ w14736;
	assign w14816 = w14741 ^ w14715;
	assign w45300 = ~w14816;
	assign w14704 = w14760 ^ w14761;
	assign w50496 = w14704 ^ w14705;
	assign w23584 = w46555 ^ w46554;
	assign w23652 = w23656 ^ w23584;
	assign w23649 = w23584 ^ w23651;
	assign w23641 = w23648 & w23652;
	assign w23573 = w23641 ^ w23570;
	assign w23577 = w23573 ^ w23571;
	assign w23582 = w46549 ^ w23577;
	assign w23545 = w23577 ^ w44360;
	assign w23588 = w46551 ^ w23545;
	assign w23640 = w23649 & w23647;
	assign w23591 = w23634 ^ w23640;
	assign w23629 = w23591 ^ w23583;
	assign w23632 = w23591 ^ w23582;
	assign w23628 = w23632 & w23631;
	assign w23623 = w23628 ^ w23588;
	assign w23622 = w23623 & w23624;
	assign w23540 = w23622 ^ w23639;
	assign w23535 = w23540 ^ w23636;
	assign w23620 = w23628 ^ w23622;
	assign w23541 = w23622 ^ w23586;
	assign w26334 = w46575 ^ w26254;
	assign w26330 = w46579 ^ w26334;
	assign w26317 = w26334 & w26330;
	assign w26222 = w26317 ^ w26266;
	assign w26304 = w46579 ^ w26222;
	assign w26270 = w26223 ^ w26224;
	assign w26269 = w26270 ^ w26252;
	assign w26311 = w26317 ^ w26269;
	assign w26308 = w26312 & w26311;
	assign w26303 = w26308 ^ w26268;
	assign w26307 = w26308 ^ w26310;
	assign w26306 = w26309 & w26307;
	assign w26217 = w26306 ^ w26318;
	assign w26213 = w26217 ^ w26253;
	assign w26212 = w46575 ^ w26213;
	assign w26214 = w26306 ^ w26262;
	assign w26305 = w26306 ^ w26268;
	assign w26275 = w26305 & w26331;
	assign w26216 = w46573 ^ w26213;
	assign w26302 = w26303 & w26304;
	assign w26221 = w26302 ^ w26266;
	assign w26301 = w26302 ^ w26310;
	assign w26300 = w26308 ^ w26302;
	assign w26220 = w26302 ^ w26319;
	assign w26287 = w26301 & w46580;
	assign w26299 = w26310 & w26300;
	assign w26297 = w26299 ^ w26307;
	assign w44470 = w26299 ^ w26317;
	assign w26291 = w44470 ^ w26269;
	assign w26280 = w26291 & w26332;
	assign w26258 = w46579 ^ w44470;
	assign w26298 = w26258 ^ w26221;
	assign w26279 = w26298 & w26329;
	assign w26296 = w26305 & w26297;
	assign w26261 = w26296 ^ w26271;
	assign w26295 = w26261 ^ w26263;
	assign w26285 = w26295 & w26334;
	assign w26292 = w26261 ^ w26214;
	assign w26219 = w26296 ^ w26320;
	assign w26211 = w26258 ^ w26219;
	assign w26290 = w26211 ^ w26212;
	assign w26282 = w26290 & w26323;
	assign w26243 = w26282 ^ w26285;
	assign w26240 = ~w26243;
	assign w26276 = w26295 & w26330;
	assign w26273 = w26290 & w26338;
	assign w26277 = w26292 & w26337;
	assign w26286 = w26292 & w26322;
	assign w26244 = w26286 ^ w26277;
	assign w26218 = w26248 ^ w26211;
	assign w44472 = w26285 ^ w26286;
	assign w26267 = w26282 ^ w44472;
	assign w26289 = w26291 & w26328;
	assign w44473 = w26287 ^ w26289;
	assign w26288 = w26298 & w26327;
	assign w26284 = w26305 & w26324;
	assign w26246 = w26284 ^ w26276;
	assign w26228 = w26284 ^ w26285;
	assign w26278 = w26301 & w26333;
	assign w26233 = w26278 ^ w26267;
	assign w26230 = ~w26233;
	assign w26215 = w26220 ^ w26316;
	assign w26294 = w26215 ^ w26218;
	assign w26272 = w26294 & w26335;
	assign w26281 = w26294 & w26326;
	assign w26259 = w26277 ^ w26281;
	assign w26237 = ~w26259;
	assign w26293 = w26215 ^ w26216;
	assign w26283 = w26293 & w26325;
	assign w26227 = w26283 ^ w26267;
	assign w26274 = w26293 & w26336;
	assign w44469 = w26273 ^ w26274;
	assign w26255 = w26279 ^ w44469;
	assign w26256 = w26280 ^ w26255;
	assign w50450 = w26256 ^ w26227;
	assign w26260 = w26288 ^ w26256;
	assign w26242 = w26246 ^ w44469;
	assign w26245 = w44473 ^ w26242;
	assign w26241 = w26237 ^ w26242;
	assign w26341 = w26240 ^ w26241;
	assign w26342 = w26244 ^ w26245;
	assign w26265 = w26289 ^ w26260;
	assign w50449 = w44472 ^ w26265;
	assign w26229 = w26287 ^ w26260;
	assign w50448 = w26228 ^ w26229;
	assign w26239 = w26282 ^ w26283;
	assign w26340 = w26265 ^ w26239;
	assign w26238 = w26283 ^ w26272;
	assign w45578 = ~w26342;
	assign w42869 = w14415 ^ w45578;
	assign w45584 = ~w26340;
	assign w45585 = ~w26341;
	assign w43054 = w45585 ^ w42876;
	assign w42873 = w45585 ^ w45289;
	assign w26234 = ~w26238;
	assign w26236 = w26237 ^ w26275;
	assign w26232 = w26236 ^ w44473;
	assign w26231 = w26255 ^ w26232;
	assign w50447 = w26230 ^ w26231;
	assign w26235 = w26274 ^ w26232;
	assign w26339 = w26234 ^ w26235;
	assign w45583 = ~w26339;
	assign w14678 = w46544 ^ w46541;
	assign w14674 = w14678 ^ w14606;
	assign w14670 = w14589 ^ w14678;
	assign w14669 = w46548 ^ w14670;
	assign w14663 = w14670 & w14674;
	assign w10844 = w46540 ^ w46534;
	assign w10914 = w10844 ^ w10839;
	assign w10924 = w46535 ^ w10844;
	assign w10920 = w46539 ^ w10924;
	assign w10907 = w10924 & w10920;
	assign w23546 = w23572 ^ w44357;
	assign w23630 = w23546 ^ w23571;
	assign w23621 = w23622 ^ w23630;
	assign w23607 = w23621 & w46556;
	assign w23627 = w23628 ^ w23630;
	assign w23626 = w23629 & w23627;
	assign w23537 = w23626 ^ w23638;
	assign w23533 = w23537 ^ w23573;
	assign w23536 = w46549 ^ w23533;
	assign w23532 = w46551 ^ w23533;
	assign w23613 = w23535 ^ w23536;
	assign w23625 = w23626 ^ w23588;
	assign w23604 = w23625 & w23644;
	assign w23534 = w23626 ^ w23582;
	assign w23603 = w23613 & w23645;
	assign w23594 = w23613 & w23656;
	assign w23598 = w23621 & w23653;
	assign w23595 = w23625 & w23651;
	assign w23619 = w23630 & w23620;
	assign w23617 = w23619 ^ w23627;
	assign w23616 = w23625 & w23617;
	assign w23539 = w23616 ^ w23640;
	assign w23581 = w23616 ^ w23591;
	assign w23615 = w23581 ^ w23583;
	assign w23612 = w23581 ^ w23534;
	assign w23605 = w23615 & w23654;
	assign w23606 = w23612 & w23642;
	assign w44361 = w23605 ^ w23606;
	assign w23597 = w23612 & w23657;
	assign w23564 = w23606 ^ w23597;
	assign w23596 = w23615 & w23650;
	assign w23566 = w23604 ^ w23596;
	assign w44359 = w23619 ^ w23637;
	assign w23578 = w46555 ^ w44359;
	assign w23618 = w23578 ^ w23541;
	assign w23599 = w23618 & w23649;
	assign w23531 = w23578 ^ w23539;
	assign w23538 = w23568 ^ w23531;
	assign w23614 = w23535 ^ w23538;
	assign w23601 = w23614 & w23646;
	assign w23610 = w23531 ^ w23532;
	assign w23602 = w23610 & w23643;
	assign w23593 = w23610 & w23658;
	assign w44358 = w23593 ^ w23594;
	assign w23575 = w23599 ^ w44358;
	assign w23562 = w23566 ^ w44358;
	assign w23579 = w23597 ^ w23601;
	assign w23592 = w23614 & w23655;
	assign w23558 = w23603 ^ w23592;
	assign w23554 = ~w23558;
	assign w23587 = w23602 ^ w44361;
	assign w23547 = w23603 ^ w23587;
	assign w23553 = w23598 ^ w23587;
	assign w23550 = ~w23553;
	assign w23608 = w23618 & w23647;
	assign w23611 = w44359 ^ w23589;
	assign w23609 = w23611 & w23648;
	assign w23600 = w23611 & w23652;
	assign w23576 = w23600 ^ w23575;
	assign w50483 = w23576 ^ w23547;
	assign w23580 = w23608 ^ w23576;
	assign w23585 = w23609 ^ w23580;
	assign w50482 = w44361 ^ w23585;
	assign w23549 = w23607 ^ w23580;
	assign w23563 = w23602 ^ w23605;
	assign w23560 = ~w23563;
	assign w23557 = ~w23579;
	assign w23561 = w23557 ^ w23562;
	assign w23661 = w23560 ^ w23561;
	assign w23556 = w23557 ^ w23595;
	assign w45507 = ~w23661;
	assign w23559 = w23602 ^ w23603;
	assign w23660 = w23585 ^ w23559;
	assign w45506 = ~w23660;
	assign w23548 = w23604 ^ w23605;
	assign w50481 = w23548 ^ w23549;
	assign w44362 = w23607 ^ w23609;
	assign w23552 = w23556 ^ w44362;
	assign w23551 = w23575 ^ w23552;
	assign w50480 = w23550 ^ w23551;
	assign w23555 = w23594 ^ w23552;
	assign w23659 = w23554 ^ w23555;
	assign w45513 = ~w23659;
	assign w23565 = w44362 ^ w23562;
	assign w23662 = w23564 ^ w23565;
	assign w45508 = ~w23662;
	assign w11365 = w11408 ^ w11409;
	assign w11466 = w11391 ^ w11365;
	assign w50292 = ~w11466;
	assign w43448 = w45313 ^ w50292;
	assign w43273 = w11466 ^ w45312;
	assign w43271 = w43272 ^ w43273;
	assign w50188 = ~w43271;
	assign w46542 = w50188 ^ w1251;
	assign w14667 = w46542 ^ w14591;
	assign w14596 = w46548 ^ w46542;
	assign w14673 = w14590 ^ w14596;
	assign w14666 = w14596 ^ w14591;
	assign w14676 = w46543 ^ w14596;
	assign w14671 = w14606 ^ w14673;
	assign w14592 = w46544 ^ w46542;
	assign w14595 = w14663 ^ w14592;
	assign w14551 = w14592 ^ w46543;
	assign w14675 = w46548 ^ w14551;
	assign w14661 = w46548 & w14675;
	assign w14672 = w46547 ^ w14676;
	assign w43257 = w43448 ^ w43419;
	assign w50197 = w50286 ^ w43257;
	assign w46533 = w50197 ^ w1260;
	assign w10926 = w46536 ^ w46533;
	assign w10905 = w10926 & w10915;
	assign w10841 = w10905 ^ w10839;
	assign w10922 = w10926 ^ w10854;
	assign w43248 = w43448 ^ w45510;
	assign w43246 = ~w43248;
	assign w50204 = w43246 ^ w43247;
	assign w46526 = w50204 ^ w1267;
	assign w26120 = w46532 ^ w46526;
	assign w26200 = w46527 ^ w26120;
	assign w26190 = w26120 ^ w26115;
	assign w26196 = w46531 ^ w26200;
	assign w26116 = w46528 ^ w46526;
	assign w26075 = w26116 ^ w46527;
	assign w26199 = w46532 ^ w26075;
	assign w26185 = w46532 & w26199;
	assign w43245 = w45321 ^ w11466;
	assign w50205 = w43244 ^ w43245;
	assign w46525 = w50205 ^ w1268;
	assign w26203 = w46525 ^ w46531;
	assign w26184 = w26203 & w26188;
	assign w43230 = w43448 ^ w43444;
	assign w50212 = w45321 ^ w43230;
	assign w46518 = w50212 ^ w1275;
	assign w29202 = w46524 ^ w46518;
	assign w29279 = w29196 ^ w29202;
	assign w26183 = w26200 & w26196;
	assign w10838 = w46535 ^ w46533;
	assign w10913 = w10838 ^ w10928;
	assign w10921 = w10838 ^ w10844;
	assign w10919 = w10854 ^ w10921;
	assign w10906 = w10921 & w10914;
	assign w10800 = w10840 ^ w10838;
	assign w10904 = w10928 & w10913;
	assign w10813 = w10904 ^ w10905;
	assign w10860 = w10813 ^ w10814;
	assign w10916 = w10837 ^ w10800;
	assign w29282 = w46519 ^ w29202;
	assign w14659 = w14676 & w14672;
	assign w10927 = w46533 ^ w46539;
	assign w10908 = w10927 & w10912;
	assign w26202 = w46528 ^ w46525;
	assign w26194 = w26113 ^ w26202;
	assign w26193 = w46532 ^ w26194;
	assign w14657 = w14678 & w14667;
	assign w14565 = w14656 ^ w14657;
	assign w14612 = w14565 ^ w14566;
	assign w14611 = w14612 ^ w14594;
	assign w14653 = w14659 ^ w14611;
	assign w10842 = w10908 ^ w10838;
	assign w10859 = w10860 ^ w10842;
	assign w10901 = w10907 ^ w10859;
	assign w26114 = w46527 ^ w46525;
	assign w26076 = w26116 ^ w26114;
	assign w26189 = w26114 ^ w26204;
	assign w26180 = w26204 & w26189;
	assign w26118 = w26184 ^ w26114;
	assign w26197 = w26114 ^ w26120;
	assign w26182 = w26197 & w26190;
	assign w26195 = w26130 ^ w26197;
	assign w26198 = w26202 ^ w26130;
	assign w26187 = w26194 & w26198;
	assign w26119 = w26187 ^ w26116;
	assign w10925 = w46533 ^ w46538;
	assign w10903 = w10925 & w10916;
	assign w43825 = w10903 ^ w10909;
	assign w10853 = w43825 ^ w10838;
	assign w43826 = w10903 ^ w10906;
	assign w10816 = w10842 ^ w43826;
	assign w10900 = w10816 ^ w10841;
	assign w10856 = w10904 ^ w43826;
	assign w10812 = w10907 ^ w10856;
	assign w14552 = w14592 ^ w14590;
	assign w14668 = w14589 ^ w14552;
	assign w14655 = w14677 & w14668;
	assign w26201 = w46525 ^ w46530;
	assign w26192 = w26113 ^ w26076;
	assign w26179 = w26201 & w26192;
	assign w44462 = w26179 ^ w26185;
	assign w26129 = w44462 ^ w26114;
	assign w44463 = w26179 ^ w26182;
	assign w26132 = w26180 ^ w44463;
	assign w26088 = w26183 ^ w26132;
	assign w26170 = w46531 ^ w26088;
	assign w26092 = w26118 ^ w44463;
	assign w14593 = w14657 ^ w14591;
	assign w14599 = w14595 ^ w14593;
	assign w14604 = w46541 ^ w14599;
	assign w26186 = w26195 & w26193;
	assign w26137 = w26180 ^ w26186;
	assign w26175 = w26137 ^ w26129;
	assign w43984 = w14655 ^ w14661;
	assign w14605 = w43984 ^ w14590;
	assign w14567 = w14599 ^ w43984;
	assign w14610 = w46543 ^ w14567;
	assign w10918 = w10837 ^ w10926;
	assign w10911 = w10918 & w10922;
	assign w10917 = w46540 ^ w10918;
	assign w10910 = w10919 & w10917;
	assign w10843 = w10911 ^ w10840;
	assign w10847 = w10843 ^ w10841;
	assign w10815 = w10847 ^ w43825;
	assign w10858 = w46535 ^ w10815;
	assign w10852 = w46533 ^ w10847;
	assign w10861 = w10904 ^ w10910;
	assign w10902 = w10861 ^ w10852;
	assign w10898 = w10902 & w10901;
	assign w10893 = w10898 ^ w10858;
	assign w10897 = w10898 ^ w10900;
	assign w10899 = w10861 ^ w10853;
	assign w10896 = w10899 & w10897;
	assign w10807 = w10896 ^ w10908;
	assign w10803 = w10807 ^ w10843;
	assign w10895 = w10896 ^ w10858;
	assign w10802 = w46535 ^ w10803;
	assign w10865 = w10895 & w10921;
	assign w10806 = w46533 ^ w10803;
	assign w10804 = w10896 ^ w10852;
	assign w10874 = w10895 & w10914;
	assign w10894 = w46539 ^ w10812;
	assign w10892 = w10893 & w10894;
	assign w10810 = w10892 ^ w10909;
	assign w10890 = w10898 ^ w10892;
	assign w10891 = w10892 ^ w10900;
	assign w10868 = w10891 & w10923;
	assign w10877 = w10891 & w46540;
	assign w10811 = w10892 ^ w10856;
	assign w10889 = w10900 & w10890;
	assign w10887 = w10889 ^ w10897;
	assign w10886 = w10895 & w10887;
	assign w10809 = w10886 ^ w10910;
	assign w10851 = w10886 ^ w10861;
	assign w10885 = w10851 ^ w10853;
	assign w10875 = w10885 & w10924;
	assign w10818 = w10874 ^ w10875;
	assign w10866 = w10885 & w10920;
	assign w10836 = w10874 ^ w10866;
	assign w10882 = w10851 ^ w10804;
	assign w10867 = w10882 & w10927;
	assign w10876 = w10882 & w10912;
	assign w10834 = w10876 ^ w10867;
	assign w43830 = w10889 ^ w10907;
	assign w10881 = w43830 ^ w10859;
	assign w10870 = w10881 & w10922;
	assign w10879 = w10881 & w10918;
	assign w43829 = w10877 ^ w10879;
	assign w10848 = w46539 ^ w43830;
	assign w10801 = w10848 ^ w10809;
	assign w10808 = w10838 ^ w10801;
	assign w10888 = w10848 ^ w10811;
	assign w10878 = w10888 & w10917;
	assign w10880 = w10801 ^ w10802;
	assign w10863 = w10880 & w10928;
	assign w10805 = w10810 ^ w10906;
	assign w10883 = w10805 ^ w10806;
	assign w10873 = w10883 & w10915;
	assign w10864 = w10883 & w10926;
	assign w43827 = w10863 ^ w10864;
	assign w10832 = w10836 ^ w43827;
	assign w10835 = w43829 ^ w10832;
	assign w10932 = w10834 ^ w10835;
	assign w10884 = w10805 ^ w10808;
	assign w10862 = w10884 & w10925;
	assign w10828 = w10873 ^ w10862;
	assign w10872 = w10880 & w10913;
	assign w10829 = w10872 ^ w10873;
	assign w10824 = ~w10828;
	assign w10833 = w10872 ^ w10875;
	assign w10830 = ~w10833;
	assign w45221 = ~w10932;
	assign w43120 = w45221 ^ w45289;
	assign w10869 = w10888 & w10919;
	assign w10845 = w10869 ^ w43827;
	assign w10846 = w10870 ^ w10845;
	assign w10850 = w10878 ^ w10846;
	assign w10819 = w10877 ^ w10850;
	assign w50452 = w10818 ^ w10819;
	assign w43144 = w50448 ^ w50452;
	assign w43026 = ~w43144;
	assign w42867 = w50459 ^ w50452;
	assign w10855 = w10879 ^ w10850;
	assign w10930 = w10855 ^ w10829;
	assign w50455 = ~w10930;
	assign w43130 = w45584 ^ w50455;
	assign w43005 = w45288 ^ w10930;
	assign w10871 = w10884 & w10916;
	assign w10849 = w10867 ^ w10871;
	assign w10827 = ~w10849;
	assign w10831 = w10827 ^ w10832;
	assign w10931 = w10830 ^ w10831;
	assign w10826 = w10827 ^ w10865;
	assign w10822 = w10826 ^ w43829;
	assign w45220 = ~w10931;
	assign w43121 = w45220 ^ w50457;
	assign w10825 = w10864 ^ w10822;
	assign w10929 = w10824 ^ w10825;
	assign w43007 = w45287 ^ w10929;
	assign w43828 = w10875 ^ w10876;
	assign w50453 = w43828 ^ w10855;
	assign w43009 = w50460 ^ w50453;
	assign w43135 = w50449 ^ w50453;
	assign w10857 = w10872 ^ w43828;
	assign w10823 = w10868 ^ w10857;
	assign w10820 = ~w10823;
	assign w50454 = ~w10929;
	assign w43132 = w45583 ^ w50454;
	assign w14658 = w14673 & w14666;
	assign w43981 = w14655 ^ w14658;
	assign w14568 = w14594 ^ w43981;
	assign w14652 = w14568 ^ w14593;
	assign w14608 = w14656 ^ w43981;
	assign w14564 = w14659 ^ w14608;
	assign w14646 = w46547 ^ w14564;
	assign w26191 = w46526 ^ w26115;
	assign w26181 = w26202 & w26191;
	assign w26089 = w26180 ^ w26181;
	assign w26117 = w26181 ^ w26115;
	assign w26123 = w26119 ^ w26117;
	assign w26128 = w46525 ^ w26123;
	assign w26176 = w26092 ^ w26117;
	assign w26136 = w26089 ^ w26090;
	assign w26178 = w26137 ^ w26128;
	assign w26091 = w26123 ^ w44462;
	assign w26134 = w46527 ^ w26091;
	assign w26135 = w26136 ^ w26118;
	assign w26177 = w26183 ^ w26135;
	assign w26174 = w26178 & w26177;
	assign w26169 = w26174 ^ w26134;
	assign w26168 = w26169 & w26170;
	assign w26166 = w26174 ^ w26168;
	assign w26167 = w26168 ^ w26176;
	assign w26144 = w26167 & w26199;
	assign w26153 = w26167 & w46532;
	assign w26087 = w26168 ^ w26132;
	assign w26086 = w26168 ^ w26185;
	assign w26165 = w26176 & w26166;
	assign w44467 = w26165 ^ w26183;
	assign w26157 = w44467 ^ w26135;
	assign w26146 = w26157 & w26198;
	assign w26124 = w46531 ^ w44467;
	assign w26164 = w26124 ^ w26087;
	assign w26145 = w26164 & w26195;
	assign w26154 = w26164 & w26193;
	assign w26081 = w26086 ^ w26182;
	assign w26173 = w26174 ^ w26176;
	assign w26163 = w26165 ^ w26173;
	assign w26172 = w26175 & w26173;
	assign w26080 = w26172 ^ w26128;
	assign w26171 = w26172 ^ w26134;
	assign w26150 = w26171 & w26190;
	assign w26141 = w26171 & w26197;
	assign w26162 = w26171 & w26163;
	assign w26127 = w26162 ^ w26137;
	assign w26158 = w26127 ^ w26080;
	assign w26143 = w26158 & w26203;
	assign w26085 = w26162 ^ w26186;
	assign w26077 = w26124 ^ w26085;
	assign w26084 = w26114 ^ w26077;
	assign w26160 = w26081 ^ w26084;
	assign w26147 = w26160 & w26192;
	assign w26138 = w26160 & w26201;
	assign w26125 = w26143 ^ w26147;
	assign w26103 = ~w26125;
	assign w26102 = w26103 ^ w26141;
	assign w26083 = w26172 ^ w26184;
	assign w26079 = w26083 ^ w26119;
	assign w26082 = w46525 ^ w26079;
	assign w26159 = w26081 ^ w26082;
	assign w26149 = w26159 & w26191;
	assign w26161 = w26127 ^ w26129;
	assign w26151 = w26161 & w26200;
	assign w26142 = w26161 & w26196;
	assign w26094 = w26150 ^ w26151;
	assign w26112 = w26150 ^ w26142;
	assign w26078 = w46527 ^ w26079;
	assign w26156 = w26077 ^ w26078;
	assign w26139 = w26156 & w26204;
	assign w26148 = w26156 & w26189;
	assign w26109 = w26148 ^ w26151;
	assign w26105 = w26148 ^ w26149;
	assign w26155 = w26157 & w26194;
	assign w44466 = w26153 ^ w26155;
	assign w26098 = w26102 ^ w44466;
	assign w26106 = ~w26109;
	assign w10817 = w10873 ^ w10857;
	assign w50456 = w10846 ^ w10817;
	assign w43080 = w50450 ^ w50456;
	assign w43081 = w50456 ^ w50461;
	assign w43015 = ~w43081;
	assign w43019 = w43015 ^ w45220;
	assign w42870 = w43080 ^ w50448;
	assign w14662 = w14671 & w14669;
	assign w14613 = w14656 ^ w14662;
	assign w14651 = w14613 ^ w14605;
	assign w14654 = w14613 ^ w14604;
	assign w14650 = w14654 & w14653;
	assign w14649 = w14650 ^ w14652;
	assign w14645 = w14650 ^ w14610;
	assign w14648 = w14651 & w14649;
	assign w14559 = w14648 ^ w14660;
	assign w14556 = w14648 ^ w14604;
	assign w14647 = w14648 ^ w14610;
	assign w14617 = w14647 & w14673;
	assign w14626 = w14647 & w14666;
	assign w14555 = w14559 ^ w14595;
	assign w14558 = w46541 ^ w14555;
	assign w14644 = w14645 & w14646;
	assign w14643 = w14644 ^ w14652;
	assign w14629 = w14643 & w46548;
	assign w14620 = w14643 & w14675;
	assign w14642 = w14650 ^ w14644;
	assign w14641 = w14652 & w14642;
	assign w14562 = w14644 ^ w14661;
	assign w14563 = w14644 ^ w14608;
	assign w43983 = w14641 ^ w14659;
	assign w14633 = w43983 ^ w14611;
	assign w14622 = w14633 & w14674;
	assign w14600 = w46547 ^ w43983;
	assign w14640 = w14600 ^ w14563;
	assign w14630 = w14640 & w14669;
	assign w14621 = w14640 & w14671;
	assign w14557 = w14562 ^ w14658;
	assign w14631 = w14633 & w14670;
	assign w43986 = w14629 ^ w14631;
	assign w14635 = w14557 ^ w14558;
	assign w14616 = w14635 & w14678;
	assign w14625 = w14635 & w14667;
	assign w14639 = w14641 ^ w14649;
	assign w14638 = w14647 & w14639;
	assign w14603 = w14638 ^ w14613;
	assign w14634 = w14603 ^ w14556;
	assign w14628 = w14634 & w14664;
	assign w14637 = w14603 ^ w14605;
	assign w14618 = w14637 & w14672;
	assign w14588 = w14626 ^ w14618;
	assign w14619 = w14634 & w14679;
	assign w14627 = w14637 & w14676;
	assign w14570 = w14626 ^ w14627;
	assign w43985 = w14627 ^ w14628;
	assign w14561 = w14638 ^ w14662;
	assign w14553 = w14600 ^ w14561;
	assign w14560 = w14590 ^ w14553;
	assign w14636 = w14557 ^ w14560;
	assign w14623 = w14636 & w14668;
	assign w14601 = w14619 ^ w14623;
	assign w14579 = ~w14601;
	assign w14614 = w14636 & w14677;
	assign w14580 = w14625 ^ w14614;
	assign w14576 = ~w14580;
	assign w14578 = w14579 ^ w14617;
	assign w14574 = w14578 ^ w43986;
	assign w14577 = w14616 ^ w14574;
	assign w14681 = w14576 ^ w14577;
	assign w45295 = ~w14681;
	assign w42987 = w45513 ^ w45295;
	assign w14554 = w46543 ^ w14555;
	assign w14632 = w14553 ^ w14554;
	assign w14624 = w14632 & w14665;
	assign w14609 = w14624 ^ w43985;
	assign w14585 = w14624 ^ w14627;
	assign w14582 = ~w14585;
	assign w14581 = w14624 ^ w14625;
	assign w14569 = w14625 ^ w14609;
	assign w14575 = w14620 ^ w14609;
	assign w14572 = ~w14575;
	assign w14615 = w14632 & w14680;
	assign w43982 = w14615 ^ w14616;
	assign w14597 = w14621 ^ w43982;
	assign w14573 = w14597 ^ w14574;
	assign w14584 = w14588 ^ w43982;
	assign w14583 = w14579 ^ w14584;
	assign w14683 = w14582 ^ w14583;
	assign w14587 = w43986 ^ w14584;
	assign w50467 = w14572 ^ w14573;
	assign w45297 = ~w14683;
	assign w26104 = w26149 ^ w26138;
	assign w26100 = ~w26104;
	assign w14598 = w14622 ^ w14597;
	assign w50470 = w14598 ^ w14569;
	assign w43086 = w50470 ^ w50483;
	assign w42837 = w43086 ^ w50481;
	assign w42833 = ~w43086;
	assign w42834 = w42833 ^ w50480;
	assign w42831 = w42833 ^ w45508;
	assign w14602 = w14630 ^ w14598;
	assign w14607 = w14631 ^ w14602;
	assign w50469 = w43985 ^ w14607;
	assign w14682 = w14607 ^ w14581;
	assign w45296 = ~w14682;
	assign w43095 = w45296 ^ w45506;
	assign w42968 = w50470 ^ w45296;
	assign w14571 = w14629 ^ w14602;
	assign w50468 = w14570 ^ w14571;
	assign w26152 = w26158 & w26188;
	assign w26110 = w26152 ^ w26143;
	assign w44465 = w26151 ^ w26152;
	assign w26133 = w26148 ^ w44465;
	assign w26093 = w26149 ^ w26133;
	assign w26099 = w26144 ^ w26133;
	assign w26096 = ~w26099;
	assign w26140 = w26159 & w26202;
	assign w44464 = w26139 ^ w26140;
	assign w26121 = w26145 ^ w44464;
	assign w26122 = w26146 ^ w26121;
	assign w50515 = w26122 ^ w26093;
	assign w26097 = w26121 ^ w26098;
	assign w50512 = w26096 ^ w26097;
	assign w26108 = w26112 ^ w44464;
	assign w26107 = w26103 ^ w26108;
	assign w26207 = w26106 ^ w26107;
	assign w26126 = w26154 ^ w26122;
	assign w26131 = w26155 ^ w26126;
	assign w26095 = w26153 ^ w26126;
	assign w50513 = w26094 ^ w26095;
	assign w26206 = w26131 ^ w26105;
	assign w50514 = w44465 ^ w26131;
	assign w42881 = w50514 ^ w50513;
	assign w26111 = w44466 ^ w26108;
	assign w26208 = w26110 ^ w26111;
	assign w45574 = ~w26208;
	assign w45580 = ~w26206;
	assign w45581 = ~w26207;
	assign w26101 = w26140 ^ w26098;
	assign w26205 = w26100 ^ w26101;
	assign w45579 = ~w26205;
	assign w43029 = w45580 ^ w45579;
	assign w14586 = w14628 ^ w14619;
	assign w14684 = w14586 ^ w14587;
	assign w45290 = ~w14684;
	assign w10821 = w10845 ^ w10822;
	assign w50451 = w10820 ^ w10821;
	assign w43119 = w50451 ^ w50458;
	assign w43002 = ~w43119;
	assign w43013 = w43144 ^ w43002;
	assign w43000 = w43002 ^ w50447;
	assign w42871 = w50447 ^ w50451;
	assign w43149 = w42870 ^ w42871;
	assign w45964 = ~w43080;
	assign w43025 = w45964 ^ w50449;
	assign w42868 = w45964 ^ w45221;
	assign w43150 = w42868 ^ w42869;
	assign w45967 = ~w43418;
	assign w43406 = w45967 ^ w45322;
	assign w43404 = w43405 ^ w43406;
	assign w50223 = ~w43404;
	assign w46507 = w50223 ^ w1223;
	assign w32769 = w46501 ^ w46507;
	assign w32762 = w46507 ^ w32766;
	assign w32696 = w46507 ^ w46506;
	assign w32749 = w32766 & w32762;
	assign w43401 = w45967 ^ w50312;
	assign w50225 = w43400 ^ w43401;
	assign w46505 = w50225 ^ w1225;
	assign w32656 = w46505 ^ w46506;
	assign w43221 = w45967 ^ w50303;
	assign w43490 = w43221 ^ w43222;
	assign w50226 = w43490 ^ w43434;
	assign w32679 = w46507 ^ w46505;
	assign w46504 = w50226 ^ w1226;
	assign w32770 = w46506 ^ w46504;
	assign w32755 = w32680 ^ w32770;
	assign w32768 = w46504 ^ w46501;
	assign w32764 = w32768 ^ w32696;
	assign w32760 = w32679 ^ w32768;
	assign w32753 = w32760 & w32764;
	assign w32746 = w32770 & w32755;
	assign w32759 = w46508 ^ w32760;
	assign w32761 = w32696 ^ w32763;
	assign w32752 = w32761 & w32759;
	assign w32703 = w32746 ^ w32752;
	assign w32681 = w46506 ^ w32679;
	assign w32756 = w32686 ^ w32681;
	assign w32748 = w32763 & w32756;
	assign w32754 = w46503 ^ w32681;
	assign w32750 = w32769 & w32754;
	assign w32684 = w32750 ^ w32680;
	assign w32757 = w46502 ^ w32681;
	assign w32747 = w32768 & w32757;
	assign w32683 = w32747 ^ w32681;
	assign w32655 = w32746 ^ w32747;
	assign w32702 = w32655 ^ w32656;
	assign w32701 = w32702 ^ w32684;
	assign w32743 = w32749 ^ w32701;
	assign w32682 = w46504 ^ w46502;
	assign w32685 = w32753 ^ w32682;
	assign w32689 = w32685 ^ w32683;
	assign w32694 = w46501 ^ w32689;
	assign w32641 = w32682 ^ w46503;
	assign w32765 = w46508 ^ w32641;
	assign w32751 = w46508 & w32765;
	assign w32642 = w32682 ^ w32680;
	assign w32744 = w32703 ^ w32694;
	assign w32740 = w32744 & w32743;
	assign w32758 = w32679 ^ w32642;
	assign w32745 = w32767 & w32758;
	assign w44738 = w32745 ^ w32751;
	assign w32657 = w32689 ^ w44738;
	assign w32695 = w44738 ^ w32680;
	assign w32741 = w32703 ^ w32695;
	assign w44739 = w32745 ^ w32748;
	assign w32698 = w32746 ^ w44739;
	assign w32654 = w32749 ^ w32698;
	assign w32658 = w32684 ^ w44739;
	assign w32742 = w32658 ^ w32683;
	assign w32739 = w32740 ^ w32742;
	assign w32738 = w32741 & w32739;
	assign w32646 = w32738 ^ w32694;
	assign w32649 = w32738 ^ w32750;
	assign w32645 = w32649 ^ w32685;
	assign w32648 = w46501 ^ w32645;
	assign w32644 = w46503 ^ w32645;
	assign w32700 = w46503 ^ w32657;
	assign w32737 = w32738 ^ w32700;
	assign w32707 = w32737 & w32763;
	assign w32735 = w32740 ^ w32700;
	assign w32716 = w32737 & w32756;
	assign w32736 = w46507 ^ w32654;
	assign w32734 = w32735 & w32736;
	assign w32652 = w32734 ^ w32751;
	assign w32647 = w32652 ^ w32748;
	assign w32725 = w32647 ^ w32648;
	assign w32706 = w32725 & w32768;
	assign w32732 = w32740 ^ w32734;
	assign w32731 = w32742 & w32732;
	assign w32733 = w32734 ^ w32742;
	assign w32653 = w32734 ^ w32698;
	assign w32715 = w32725 & w32757;
	assign w32710 = w32733 & w32765;
	assign w32719 = w32733 & w46508;
	assign w44743 = w32731 ^ w32749;
	assign w32690 = w46507 ^ w44743;
	assign w32730 = w32690 ^ w32653;
	assign w32711 = w32730 & w32761;
	assign w32720 = w32730 & w32759;
	assign w32723 = w44743 ^ w32701;
	assign w32721 = w32723 & w32760;
	assign w44742 = w32719 ^ w32721;
	assign w32712 = w32723 & w32764;
	assign w32729 = w32731 ^ w32739;
	assign w32728 = w32737 & w32729;
	assign w32651 = w32728 ^ w32752;
	assign w32643 = w32690 ^ w32651;
	assign w32722 = w32643 ^ w32644;
	assign w32714 = w32722 & w32755;
	assign w32650 = w32680 ^ w32643;
	assign w32726 = w32647 ^ w32650;
	assign w32704 = w32726 & w32767;
	assign w32693 = w32728 ^ w32703;
	assign w32724 = w32693 ^ w32646;
	assign w32709 = w32724 & w32769;
	assign w32713 = w32726 & w32758;
	assign w32691 = w32709 ^ w32713;
	assign w32669 = ~w32691;
	assign w32668 = w32669 ^ w32707;
	assign w32664 = w32668 ^ w44742;
	assign w32667 = w32706 ^ w32664;
	assign w32671 = w32714 ^ w32715;
	assign w32718 = w32724 & w32754;
	assign w32676 = w32718 ^ w32709;
	assign w32727 = w32693 ^ w32695;
	assign w32708 = w32727 & w32762;
	assign w32678 = w32716 ^ w32708;
	assign w32717 = w32727 & w32766;
	assign w32660 = w32716 ^ w32717;
	assign w32675 = w32714 ^ w32717;
	assign w32672 = ~w32675;
	assign w44741 = w32717 ^ w32718;
	assign w32699 = w32714 ^ w44741;
	assign w32665 = w32710 ^ w32699;
	assign w32662 = ~w32665;
	assign w32659 = w32715 ^ w32699;
	assign w32705 = w32722 & w32770;
	assign w44740 = w32705 ^ w32706;
	assign w32687 = w32711 ^ w44740;
	assign w32663 = w32687 ^ w32664;
	assign w32688 = w32712 ^ w32687;
	assign w50475 = w32688 ^ w32659;
	assign w43077 = w50470 ^ w50475;
	assign w42940 = w43077 ^ w45506;
	assign w32692 = w32720 ^ w32688;
	assign w32661 = w32719 ^ w32692;
	assign w50473 = w32660 ^ w32661;
	assign w43109 = w50468 ^ w50473;
	assign w42973 = ~w43109;
	assign w42836 = ~w50473;
	assign w42835 = w42836 ^ w50467;
	assign w43164 = w42834 ^ w42835;
	assign w32697 = w32721 ^ w32692;
	assign w50474 = w44741 ^ w32697;
	assign w42838 = w50474 ^ w50468;
	assign w43105 = w50469 ^ w50474;
	assign w42947 = ~w43105;
	assign w43163 = w42837 ^ w42838;
	assign w32772 = w32697 ^ w32671;
	assign w32674 = w32678 ^ w44740;
	assign w32677 = w44742 ^ w32674;
	assign w32774 = w32676 ^ w32677;
	assign w32673 = w32669 ^ w32674;
	assign w32773 = w32672 ^ w32673;
	assign w50471 = ~w32773;
	assign w43116 = w45297 ^ w50471;
	assign w42832 = w32773 ^ w45290;
	assign w43165 = w42831 ^ w42832;
	assign w50472 = w32662 ^ w32663;
	assign w43112 = w50467 ^ w50472;
	assign w42991 = w50472 ^ w45297;
	assign w42965 = ~w43112;
	assign w42963 = w42965 ^ w50480;
	assign w45758 = ~w32774;
	assign w43117 = w45290 ^ w45758;
	assign w45765 = ~w32772;
	assign w32670 = w32715 ^ w32704;
	assign w32666 = ~w32670;
	assign w32771 = w32666 ^ w32667;
	assign w45764 = ~w32771;
	assign w43101 = w45295 ^ w45764;
	assign w42989 = w45764 ^ w50469;
	assign w42969 = w43101 ^ w43095;
	assign w42962 = w43101 ^ w45513;
	assign w42960 = ~w42962;
	assign w42959 = w45765 ^ w45764;
	assign w45966 = ~w43077;
	assign w42979 = w45966 ^ w45297;
	assign w42975 = w45966 ^ w50468;
	assign w42972 = w45966 ^ w50469;
	assign w45968 = ~w43417;
	assign w43408 = w45968 ^ w45670;
	assign w50221 = w43408 ^ w43409;
	assign w43380 = w45968 ^ w45310;
	assign w50239 = w43379 ^ w43380;
	assign w46491 = w50239 ^ w1239;
	assign w29151 = w46485 ^ w46491;
	assign w29078 = w46491 ^ w46490;
	assign w29143 = w29078 ^ w29145;
	assign w29146 = w29150 ^ w29078;
	assign w29144 = w46491 ^ w29148;
	assign w29131 = w29148 & w29144;
	assign w43377 = w45968 ^ w50303;
	assign w43375 = w43376 ^ w43377;
	assign w50241 = ~w43375;
	assign w46489 = w50241 ^ w1241;
	assign w29061 = w46491 ^ w46489;
	assign w29063 = w46490 ^ w29061;
	assign w29136 = w46487 ^ w29063;
	assign w29139 = w46486 ^ w29063;
	assign w29138 = w29068 ^ w29063;
	assign w29142 = w29061 ^ w29150;
	assign w29135 = w29142 & w29146;
	assign w29132 = w29151 & w29136;
	assign w29066 = w29132 ^ w29062;
	assign w29130 = w29145 & w29138;
	assign w29129 = w29150 & w29139;
	assign w29037 = w29128 ^ w29129;
	assign w29065 = w29129 ^ w29063;
	assign w29140 = w29061 ^ w29024;
	assign w29127 = w29149 & w29140;
	assign w29067 = w29135 ^ w29064;
	assign w29071 = w29067 ^ w29065;
	assign w29076 = w46485 ^ w29071;
	assign w29141 = w46492 ^ w29142;
	assign w29134 = w29143 & w29141;
	assign w29085 = w29128 ^ w29134;
	assign w29038 = w46489 ^ w46490;
	assign w29084 = w29037 ^ w29038;
	assign w29083 = w29084 ^ w29066;
	assign w29125 = w29131 ^ w29083;
	assign w44586 = w29127 ^ w29133;
	assign w29039 = w29071 ^ w44586;
	assign w29082 = w46487 ^ w29039;
	assign w29077 = w44586 ^ w29062;
	assign w29123 = w29085 ^ w29077;
	assign w44587 = w29127 ^ w29130;
	assign w29080 = w29128 ^ w44587;
	assign w29036 = w29131 ^ w29080;
	assign w29118 = w46491 ^ w29036;
	assign w46509 = w50221 ^ w1221;
	assign w14543 = w46509 ^ w46514;
	assign w14456 = w46511 ^ w46509;
	assign w14539 = w14456 ^ w14462;
	assign w14537 = w14472 ^ w14539;
	assign w14544 = w46512 ^ w46509;
	assign w14536 = w14455 ^ w14544;
	assign w14545 = w46509 ^ w46515;
	assign w14540 = w14544 ^ w14472;
	assign w14529 = w14536 & w14540;
	assign w14461 = w14529 ^ w14458;
	assign w14523 = w14544 & w14533;
	assign w14459 = w14523 ^ w14457;
	assign w14465 = w14461 ^ w14459;
	assign w14470 = w46509 ^ w14465;
	assign w14526 = w14545 & w14530;
	assign w14460 = w14526 ^ w14456;
	assign w14418 = w14458 ^ w14456;
	assign w14534 = w14455 ^ w14418;
	assign w14521 = w14543 & w14534;
	assign w43975 = w14521 ^ w14527;
	assign w14433 = w14465 ^ w43975;
	assign w14476 = w46511 ^ w14433;
	assign w14471 = w43975 ^ w14456;
	assign w14535 = w46516 ^ w14536;
	assign w14528 = w14537 & w14535;
	assign w14524 = w14539 & w14532;
	assign w43976 = w14521 ^ w14524;
	assign w14434 = w14460 ^ w43976;
	assign w14518 = w14434 ^ w14459;
	assign w29040 = w29066 ^ w44587;
	assign w29124 = w29040 ^ w29065;
	assign w14531 = w14456 ^ w14546;
	assign w14522 = w14546 & w14531;
	assign w14474 = w14522 ^ w43976;
	assign w14430 = w14525 ^ w14474;
	assign w14431 = w14522 ^ w14523;
	assign w14512 = w46515 ^ w14430;
	assign w14479 = w14522 ^ w14528;
	assign w14520 = w14479 ^ w14470;
	assign w14517 = w14479 ^ w14471;
	assign w29126 = w29085 ^ w29076;
	assign w29122 = w29126 & w29125;
	assign w29121 = w29122 ^ w29124;
	assign w29117 = w29122 ^ w29082;
	assign w29116 = w29117 & w29118;
	assign w29034 = w29116 ^ w29133;
	assign w29114 = w29122 ^ w29116;
	assign w29113 = w29124 & w29114;
	assign w29115 = w29116 ^ w29124;
	assign w29101 = w29115 & w46492;
	assign w29092 = w29115 & w29147;
	assign w29111 = w29113 ^ w29121;
	assign w29035 = w29116 ^ w29080;
	assign w29029 = w29034 ^ w29130;
	assign w44591 = w29113 ^ w29131;
	assign w29105 = w44591 ^ w29083;
	assign w29094 = w29105 & w29146;
	assign w29103 = w29105 & w29142;
	assign w44590 = w29101 ^ w29103;
	assign w29072 = w46491 ^ w44591;
	assign w29112 = w29072 ^ w29035;
	assign w29102 = w29112 & w29141;
	assign w29093 = w29112 & w29143;
	assign w29120 = w29123 & w29121;
	assign w29028 = w29120 ^ w29076;
	assign w29031 = w29120 ^ w29132;
	assign w29027 = w29031 ^ w29067;
	assign w29119 = w29120 ^ w29082;
	assign w29110 = w29119 & w29111;
	assign w29075 = w29110 ^ w29085;
	assign w29106 = w29075 ^ w29028;
	assign w29109 = w29075 ^ w29077;
	assign w29099 = w29109 & w29148;
	assign w29098 = w29119 & w29138;
	assign w29091 = w29106 & w29151;
	assign w29090 = w29109 & w29144;
	assign w29089 = w29119 & w29145;
	assign w29100 = w29106 & w29136;
	assign w29058 = w29100 ^ w29091;
	assign w29033 = w29110 ^ w29134;
	assign w29025 = w29072 ^ w29033;
	assign w29032 = w29062 ^ w29025;
	assign w29108 = w29029 ^ w29032;
	assign w29095 = w29108 & w29140;
	assign w29073 = w29091 ^ w29095;
	assign w29086 = w29108 & w29149;
	assign w29026 = w46487 ^ w29027;
	assign w29104 = w29025 ^ w29026;
	assign w29096 = w29104 & w29137;
	assign w29087 = w29104 & w29152;
	assign w44589 = w29099 ^ w29100;
	assign w29081 = w29096 ^ w44589;
	assign w29047 = w29092 ^ w29081;
	assign w29044 = ~w29047;
	assign w29051 = ~w29073;
	assign w29050 = w29051 ^ w29089;
	assign w29046 = w29050 ^ w44590;
	assign w29057 = w29096 ^ w29099;
	assign w29054 = ~w29057;
	assign w29060 = w29098 ^ w29090;
	assign w29030 = w46485 ^ w29027;
	assign w29107 = w29029 ^ w29030;
	assign w29088 = w29107 & w29150;
	assign w29097 = w29107 & w29139;
	assign w29049 = w29088 ^ w29046;
	assign w44588 = w29087 ^ w29088;
	assign w29069 = w29093 ^ w44588;
	assign w29070 = w29094 ^ w29069;
	assign w29074 = w29102 ^ w29070;
	assign w29043 = w29101 ^ w29074;
	assign w29079 = w29103 ^ w29074;
	assign w50518 = w44589 ^ w29079;
	assign w43090 = w50514 ^ w50518;
	assign w29041 = w29097 ^ w29081;
	assign w50519 = w29070 ^ w29041;
	assign w43073 = w50515 ^ w50519;
	assign w29052 = w29097 ^ w29086;
	assign w29048 = ~w29052;
	assign w29153 = w29048 ^ w29049;
	assign w29045 = w29069 ^ w29046;
	assign w50516 = w29044 ^ w29045;
	assign w43091 = w50512 ^ w50516;
	assign w29056 = w29060 ^ w44588;
	assign w29055 = w29051 ^ w29056;
	assign w29155 = w29054 ^ w29055;
	assign w45658 = ~w29155;
	assign w43103 = w45581 ^ w45658;
	assign w45664 = ~w29153;
	assign w29059 = w44590 ^ w29056;
	assign w29156 = w29058 ^ w29059;
	assign w45659 = ~w29156;
	assign w43123 = w45574 ^ w45659;
	assign w29053 = w29096 ^ w29097;
	assign w29154 = w29079 ^ w29053;
	assign w45665 = ~w29154;
	assign w43096 = w45580 ^ w45665;
	assign w29042 = w29098 ^ w29099;
	assign w50517 = w29042 ^ w29043;
	assign w42880 = w43073 ^ w50517;
	assign w43145 = w42880 ^ w42881;
	assign w42842 = w50517 ^ w50516;
	assign w45963 = ~w43073;
	assign w43064 = w45963 ^ w45665;
	assign w43036 = w45963 ^ w45581;
	assign w14478 = w14431 ^ w14432;
	assign w14477 = w14478 ^ w14460;
	assign w14519 = w14525 ^ w14477;
	assign w14516 = w14520 & w14519;
	assign w14515 = w14516 ^ w14518;
	assign w14514 = w14517 & w14515;
	assign w14425 = w14514 ^ w14526;
	assign w14421 = w14425 ^ w14461;
	assign w14424 = w46509 ^ w14421;
	assign w14511 = w14516 ^ w14476;
	assign w14510 = w14511 & w14512;
	assign w14509 = w14510 ^ w14518;
	assign w14486 = w14509 & w14541;
	assign w14428 = w14510 ^ w14527;
	assign w14423 = w14428 ^ w14524;
	assign w14501 = w14423 ^ w14424;
	assign w14482 = w14501 & w14544;
	assign w14491 = w14501 & w14533;
	assign w14429 = w14510 ^ w14474;
	assign w14422 = w14514 ^ w14470;
	assign w14420 = w46511 ^ w14421;
	assign w14508 = w14516 ^ w14510;
	assign w14507 = w14518 & w14508;
	assign w14505 = w14507 ^ w14515;
	assign w43980 = w14507 ^ w14525;
	assign w14499 = w43980 ^ w14477;
	assign w14466 = w46515 ^ w43980;
	assign w14506 = w14466 ^ w14429;
	assign w14487 = w14506 & w14537;
	assign w14495 = w14509 & w46516;
	assign w14488 = w14499 & w14540;
	assign w14513 = w14514 ^ w14476;
	assign w14483 = w14513 & w14539;
	assign w14492 = w14513 & w14532;
	assign w14504 = w14513 & w14505;
	assign w14427 = w14504 ^ w14528;
	assign w14419 = w14466 ^ w14427;
	assign w14426 = w14456 ^ w14419;
	assign w14502 = w14423 ^ w14426;
	assign w14480 = w14502 & w14543;
	assign w14498 = w14419 ^ w14420;
	assign w14481 = w14498 & w14546;
	assign w14490 = w14498 & w14531;
	assign w14447 = w14490 ^ w14491;
	assign w14489 = w14502 & w14534;
	assign w43977 = w14481 ^ w14482;
	assign w14463 = w14487 ^ w43977;
	assign w14464 = w14488 ^ w14463;
	assign w14469 = w14504 ^ w14479;
	assign w14503 = w14469 ^ w14471;
	assign w14484 = w14503 & w14538;
	assign w14454 = w14492 ^ w14484;
	assign w14450 = w14454 ^ w43977;
	assign w14493 = w14503 & w14542;
	assign w14451 = w14490 ^ w14493;
	assign w14448 = ~w14451;
	assign w14436 = w14492 ^ w14493;
	assign w14500 = w14469 ^ w14422;
	assign w14485 = w14500 & w14545;
	assign w14494 = w14500 & w14530;
	assign w14452 = w14494 ^ w14485;
	assign w43978 = w14493 ^ w14494;
	assign w14475 = w14490 ^ w43978;
	assign w14435 = w14491 ^ w14475;
	assign w50487 = w14464 ^ w14435;
	assign w14441 = w14486 ^ w14475;
	assign w14438 = ~w14441;
	assign w14496 = w14506 & w14535;
	assign w14468 = w14496 ^ w14464;
	assign w14437 = w14495 ^ w14468;
	assign w50485 = w14436 ^ w14437;
	assign w14467 = w14485 ^ w14489;
	assign w14445 = ~w14467;
	assign w14444 = w14445 ^ w14483;
	assign w14449 = w14445 ^ w14450;
	assign w14549 = w14448 ^ w14449;
	assign w45293 = ~w14549;
	assign w14497 = w14499 & w14536;
	assign w14473 = w14497 ^ w14468;
	assign w50486 = w43978 ^ w14473;
	assign w14548 = w14473 ^ w14447;
	assign w43979 = w14495 ^ w14497;
	assign w14453 = w43979 ^ w14450;
	assign w14550 = w14452 ^ w14453;
	assign w14440 = w14444 ^ w43979;
	assign w14443 = w14482 ^ w14440;
	assign w14439 = w14463 ^ w14440;
	assign w50484 = w14438 ^ w14439;
	assign w45286 = ~w14550;
	assign w45292 = ~w14548;
	assign w14446 = w14491 ^ w14480;
	assign w14442 = ~w14446;
	assign w14547 = w14442 ^ w14443;
	assign w45291 = ~w14547;
	assign w45969 = ~w43424;
	assign w43369 = w45969 ^ w50248;
	assign w50130 = w43368 ^ w43369;
	assign w46600 = w50130 ^ w1321;
	assign w32902 = w46600 ^ w46597;
	assign w32904 = w46602 ^ w46600;
	assign w32889 = w32814 ^ w32904;
	assign w32816 = w46600 ^ w46598;
	assign w32776 = w32816 ^ w32814;
	assign w32880 = w32904 & w32889;
	assign w43348 = w45969 ^ w50265;
	assign w50141 = w43348 ^ w43349;
	assign w46589 = w50141 ^ w1332;
	assign w14946 = w46592 ^ w46589;
	assign w14925 = w14946 & w14935;
	assign w14858 = w46591 ^ w46589;
	assign w14933 = w14858 ^ w14948;
	assign w14941 = w14858 ^ w14864;
	assign w14942 = w14946 ^ w14874;
	assign w14924 = w14948 & w14933;
	assign w14833 = w14924 ^ w14925;
	assign w14880 = w14833 ^ w14834;
	assign w14938 = w14857 ^ w14946;
	assign w14931 = w14938 & w14942;
	assign w43212 = w45969 ^ w45228;
	assign w43494 = w43212 ^ w43213;
	assign w50127 = w43494 ^ w43486;
	assign w46603 = w50127 ^ w1318;
	assign w32813 = w46603 ^ w46601;
	assign w32815 = w46602 ^ w32813;
	assign w32890 = w32820 ^ w32815;
	assign w32882 = w32897 & w32890;
	assign w32896 = w46603 ^ w32900;
	assign w32883 = w32900 & w32896;
	assign w32830 = w46603 ^ w46602;
	assign w32898 = w32902 ^ w32830;
	assign w32895 = w32830 ^ w32897;
	assign w32891 = w46598 ^ w32815;
	assign w32881 = w32902 & w32891;
	assign w32817 = w32881 ^ w32815;
	assign w32903 = w46597 ^ w46603;
	assign w14937 = w46596 ^ w14938;
	assign w14863 = w14931 ^ w14860;
	assign w14861 = w14925 ^ w14859;
	assign w14867 = w14863 ^ w14861;
	assign w14872 = w46589 ^ w14867;
	assign w32894 = w32813 ^ w32902;
	assign w32893 = w46604 ^ w32894;
	assign w32886 = w32895 & w32893;
	assign w32887 = w32894 & w32898;
	assign w32819 = w32887 ^ w32816;
	assign w32823 = w32819 ^ w32817;
	assign w32828 = w46597 ^ w32823;
	assign w14939 = w14874 ^ w14941;
	assign w14930 = w14939 & w14937;
	assign w14926 = w14941 & w14934;
	assign w14820 = w14860 ^ w14858;
	assign w14936 = w14857 ^ w14820;
	assign w14881 = w14924 ^ w14930;
	assign w14922 = w14881 ^ w14872;
	assign w14947 = w46589 ^ w46595;
	assign w14928 = w14947 & w14932;
	assign w14862 = w14928 ^ w14858;
	assign w14879 = w14880 ^ w14862;
	assign w14921 = w14927 ^ w14879;
	assign w14918 = w14922 & w14921;
	assign w32892 = w32813 ^ w32776;
	assign w32879 = w32901 & w32892;
	assign w44745 = w32879 ^ w32882;
	assign w32832 = w32880 ^ w44745;
	assign w32788 = w32883 ^ w32832;
	assign w32870 = w46603 ^ w32788;
	assign w32789 = w32880 ^ w32881;
	assign w32836 = w32789 ^ w32790;
	assign w32775 = w32816 ^ w46599;
	assign w32899 = w46604 ^ w32775;
	assign w32885 = w46604 & w32899;
	assign w44744 = w32879 ^ w32885;
	assign w32829 = w44744 ^ w32814;
	assign w32791 = w32823 ^ w44744;
	assign w32834 = w46599 ^ w32791;
	assign w32837 = w32880 ^ w32886;
	assign w32878 = w32837 ^ w32828;
	assign w32875 = w32837 ^ w32829;
	assign w32888 = w46599 ^ w32815;
	assign w32884 = w32903 & w32888;
	assign w32818 = w32884 ^ w32814;
	assign w32792 = w32818 ^ w44745;
	assign w32835 = w32836 ^ w32818;
	assign w32877 = w32883 ^ w32835;
	assign w32874 = w32878 & w32877;
	assign w32869 = w32874 ^ w32834;
	assign w32868 = w32869 & w32870;
	assign w32787 = w32868 ^ w32832;
	assign w32866 = w32874 ^ w32868;
	assign w32876 = w32792 ^ w32817;
	assign w32867 = w32868 ^ w32876;
	assign w32844 = w32867 & w32899;
	assign w32873 = w32874 ^ w32876;
	assign w32872 = w32875 & w32873;
	assign w32871 = w32872 ^ w32834;
	assign w32865 = w32876 & w32866;
	assign w32863 = w32865 ^ w32873;
	assign w32841 = w32871 & w32897;
	assign w32850 = w32871 & w32890;
	assign w32853 = w32867 & w46604;
	assign w44748 = w32865 ^ w32883;
	assign w32857 = w44748 ^ w32835;
	assign w32855 = w32857 & w32894;
	assign w32846 = w32857 & w32898;
	assign w44747 = w32853 ^ w32855;
	assign w32824 = w46603 ^ w44748;
	assign w32864 = w32824 ^ w32787;
	assign w32845 = w32864 & w32895;
	assign w32862 = w32871 & w32863;
	assign w32827 = w32862 ^ w32837;
	assign w32861 = w32827 ^ w32829;
	assign w32842 = w32861 & w32896;
	assign w32812 = w32850 ^ w32842;
	assign w32851 = w32861 & w32900;
	assign w32794 = w32850 ^ w32851;
	assign w32785 = w32862 ^ w32886;
	assign w32777 = w32824 ^ w32785;
	assign w32784 = w32814 ^ w32777;
	assign w32854 = w32864 & w32893;
	assign w32783 = w32872 ^ w32884;
	assign w32779 = w32783 ^ w32819;
	assign w32782 = w46597 ^ w32779;
	assign w32778 = w46599 ^ w32779;
	assign w32856 = w32777 ^ w32778;
	assign w32839 = w32856 & w32904;
	assign w32780 = w32872 ^ w32828;
	assign w32858 = w32827 ^ w32780;
	assign w32843 = w32858 & w32903;
	assign w32852 = w32858 & w32888;
	assign w32810 = w32852 ^ w32843;
	assign w44746 = w32851 ^ w32852;
	assign w32848 = w32856 & w32889;
	assign w32833 = w32848 ^ w44746;
	assign w32809 = w32848 ^ w32851;
	assign w32806 = ~w32809;
	assign w32799 = w32844 ^ w32833;
	assign w32796 = ~w32799;
	assign w14945 = w46589 ^ w46594;
	assign w14923 = w14945 & w14936;
	assign w43993 = w14923 ^ w14926;
	assign w14876 = w14924 ^ w43993;
	assign w14832 = w14927 ^ w14876;
	assign w14914 = w46595 ^ w14832;
	assign w43992 = w14923 ^ w14929;
	assign w14835 = w14867 ^ w43992;
	assign w14878 = w46591 ^ w14835;
	assign w14873 = w43992 ^ w14858;
	assign w14913 = w14918 ^ w14878;
	assign w14912 = w14913 & w14914;
	assign w14910 = w14918 ^ w14912;
	assign w14830 = w14912 ^ w14929;
	assign w14825 = w14830 ^ w14926;
	assign w14919 = w14881 ^ w14873;
	assign w14836 = w14862 ^ w43993;
	assign w14831 = w14912 ^ w14876;
	assign w14920 = w14836 ^ w14861;
	assign w14917 = w14918 ^ w14920;
	assign w14916 = w14919 & w14917;
	assign w14827 = w14916 ^ w14928;
	assign w14824 = w14916 ^ w14872;
	assign w14823 = w14827 ^ w14863;
	assign w14822 = w46591 ^ w14823;
	assign w14826 = w46589 ^ w14823;
	assign w14903 = w14825 ^ w14826;
	assign w14915 = w14916 ^ w14878;
	assign w14885 = w14915 & w14941;
	assign w14911 = w14912 ^ w14920;
	assign w14897 = w14911 & w46596;
	assign w14888 = w14911 & w14943;
	assign w14894 = w14915 & w14934;
	assign w14893 = w14903 & w14935;
	assign w14909 = w14920 & w14910;
	assign w14907 = w14909 ^ w14917;
	assign w14906 = w14915 & w14907;
	assign w14871 = w14906 ^ w14881;
	assign w14902 = w14871 ^ w14824;
	assign w14887 = w14902 & w14947;
	assign w14896 = w14902 & w14932;
	assign w43996 = w14909 ^ w14927;
	assign w14868 = w46595 ^ w43996;
	assign w14901 = w43996 ^ w14879;
	assign w14899 = w14901 & w14938;
	assign w14890 = w14901 & w14942;
	assign w43995 = w14897 ^ w14899;
	assign w14905 = w14871 ^ w14873;
	assign w14895 = w14905 & w14944;
	assign w14838 = w14894 ^ w14895;
	assign w14886 = w14905 & w14940;
	assign w43994 = w14895 ^ w14896;
	assign w14854 = w14896 ^ w14887;
	assign w14908 = w14868 ^ w14831;
	assign w14898 = w14908 & w14937;
	assign w14829 = w14906 ^ w14930;
	assign w14821 = w14868 ^ w14829;
	assign w14828 = w14858 ^ w14821;
	assign w14900 = w14821 ^ w14822;
	assign w14904 = w14825 ^ w14828;
	assign w14891 = w14904 & w14936;
	assign w14869 = w14887 ^ w14891;
	assign w14882 = w14904 & w14945;
	assign w14848 = w14893 ^ w14882;
	assign w14847 = ~w14869;
	assign w14844 = ~w14848;
	assign w14892 = w14900 & w14933;
	assign w14853 = w14892 ^ w14895;
	assign w14877 = w14892 ^ w43994;
	assign w14837 = w14893 ^ w14877;
	assign w14849 = w14892 ^ w14893;
	assign w14883 = w14900 & w14948;
	assign w14889 = w14908 & w14939;
	assign w14884 = w14903 & w14946;
	assign w14846 = w14847 ^ w14885;
	assign w14856 = w14894 ^ w14886;
	assign w43539 = w14883 ^ w14884;
	assign w14865 = w14889 ^ w43539;
	assign w14866 = w14890 ^ w14865;
	assign w50479 = w14866 ^ w14837;
	assign w43076 = w50479 ^ w50483;
	assign w43084 = w50475 ^ w50479;
	assign w42985 = w43095 ^ w43076;
	assign w50358 = w50475 ^ w42985;
	assign w42967 = w43076 ^ w45765;
	assign w50366 = w42967 ^ w42968;
	assign w46437 = w50366 ^ w431;
	assign w42966 = w43117 ^ w43084;
	assign w50367 = w45508 ^ w42966;
	assign w46436 = w50367 ^ w432;
	assign w42956 = w43117 ^ w43076;
	assign w42849 = ~w43084;
	assign w42847 = w42849 ^ w50482;
	assign w42845 = w43084 ^ w50481;
	assign w42843 = w43084 ^ w45507;
	assign w46445 = w50358 ^ w423;
	assign w14870 = w14898 ^ w14866;
	assign w14839 = w14897 ^ w14870;
	assign w50477 = w14838 ^ w14839;
	assign w43102 = w50477 ^ w50481;
	assign w42952 = w43076 ^ w50477;
	assign w50354 = w43164 ^ w43102;
	assign w46449 = w50354 ^ w419;
	assign w42974 = w42965 ^ w43102;
	assign w50362 = w42974 ^ w42975;
	assign w46441 = w50362 ^ w427;
	assign w42944 = w42947 ^ w43102;
	assign w14875 = w14899 ^ w14870;
	assign w14950 = w14875 ^ w14849;
	assign w45304 = ~w14950;
	assign w43094 = w45765 ^ w45304;
	assign w42986 = w43094 ^ w45506;
	assign w50357 = w42986 ^ w42987;
	assign w50365 = w45304 ^ w42969;
	assign w46438 = w50365 ^ w430;
	assign w42957 = w43094 ^ w43077;
	assign w50374 = w50483 ^ w42957;
	assign w46429 = w50374 ^ w439;
	assign w42941 = w50479 ^ w45304;
	assign w50382 = w42940 ^ w42941;
	assign w46421 = w50382 ^ w447;
	assign w46446 = w50357 ^ w422;
	assign w50478 = w43994 ^ w14875;
	assign w43097 = w50478 ^ w50482;
	assign w42943 = w43101 ^ w43097;
	assign w50355 = w43163 ^ w43097;
	assign w46448 = w50355 ^ w420;
	assign w14142 = w46448 ^ w46445;
	assign w42971 = w42973 ^ w43097;
	assign w50363 = w42971 ^ w42972;
	assign w46440 = w50363 ^ w428;
	assign w10572 = w46440 ^ w46438;
	assign w10658 = w46440 ^ w46437;
	assign w42946 = ~w50478;
	assign w42961 = w42946 ^ w50474;
	assign w42945 = w43076 ^ w42946;
	assign w50379 = w42944 ^ w42945;
	assign w46424 = w50379 ^ w444;
	assign w39602 = w46424 ^ w46421;
	assign w14056 = w46448 ^ w46446;
	assign w50372 = w42960 ^ w42961;
	assign w42848 = w50477 ^ w42836;
	assign w43158 = w42847 ^ w42848;
	assign w50371 = w43158 ^ w43105;
	assign w46432 = w50371 ^ w436;
	assign w40272 = w46432 ^ w46429;
	assign w14852 = w14856 ^ w43539;
	assign w14851 = w14847 ^ w14852;
	assign w14855 = w43995 ^ w14852;
	assign w14952 = w14854 ^ w14855;
	assign w45298 = ~w14952;
	assign w43114 = w45298 ^ w45508;
	assign w42992 = w43114 ^ w43086;
	assign w50351 = w45758 ^ w42992;
	assign w46452 = w50351 ^ w416;
	assign w14060 = w46452 ^ w46446;
	assign w42980 = w43114 ^ w43077;
	assign w50359 = w45290 ^ w42980;
	assign w50375 = w45298 ^ w42956;
	assign w42954 = w43116 ^ w43114;
	assign w42844 = w45298 ^ w45758;
	assign w43160 = w42843 ^ w42844;
	assign w50368 = w43160 ^ w43116;
	assign w46435 = w50368 ^ w433;
	assign w40273 = w46429 ^ w46435;
	assign w46444 = w50359 ^ w424;
	assign w10576 = w46444 ^ w46438;
	assign w46428 = w50375 ^ w440;
	assign w14842 = w14846 ^ w43995;
	assign w14841 = w14865 ^ w14842;
	assign w14845 = w14884 ^ w14842;
	assign w14949 = w14844 ^ w14845;
	assign w45303 = ~w14949;
	assign w43092 = w45303 ^ w45513;
	assign w42988 = w43092 ^ w50482;
	assign w50356 = w42988 ^ w42989;
	assign w42970 = w43105 ^ w43092;
	assign w50364 = w45295 ^ w42970;
	assign w42958 = w43095 ^ w45303;
	assign w50373 = w42958 ^ w42959;
	assign w50380 = w45303 ^ w42943;
	assign w46423 = w50380 ^ w445;
	assign w39514 = w46423 ^ w46421;
	assign w42942 = w43094 ^ w43092;
	assign w50381 = w45296 ^ w42942;
	assign w46422 = w50381 ^ w446;
	assign w39516 = w46424 ^ w46422;
	assign w39520 = w46428 ^ w46422;
	assign w39597 = w39514 ^ w39520;
	assign w39600 = w46423 ^ w39520;
	assign w39476 = w39516 ^ w39514;
	assign w39475 = w39516 ^ w46423;
	assign w39599 = w46428 ^ w39475;
	assign w39585 = w46428 & w39599;
	assign w46430 = w50373 ^ w438;
	assign w40186 = w46432 ^ w46430;
	assign w40190 = w46436 ^ w46430;
	assign w46447 = w50356 ^ w421;
	assign w14054 = w46447 ^ w46445;
	assign w14137 = w14054 ^ w14060;
	assign w14015 = w14056 ^ w46447;
	assign w14140 = w46447 ^ w14060;
	assign w46439 = w50364 ^ w429;
	assign w10656 = w46439 ^ w10576;
	assign w10531 = w10572 ^ w46439;
	assign w10655 = w46444 ^ w10531;
	assign w10641 = w46444 & w10655;
	assign w14016 = w14056 ^ w14054;
	assign w14139 = w46452 ^ w14015;
	assign w14125 = w46452 & w14139;
	assign w10570 = w46439 ^ w46437;
	assign w10653 = w10570 ^ w10576;
	assign w10532 = w10572 ^ w10570;
	assign w46431 = w50372 ^ w437;
	assign w40184 = w46431 ^ w46429;
	assign w40267 = w40184 ^ w40190;
	assign w40270 = w46431 ^ w40190;
	assign w40266 = w46435 ^ w40270;
	assign w40146 = w40186 ^ w40184;
	assign w40145 = w40186 ^ w46431;
	assign w40269 = w46436 ^ w40145;
	assign w40255 = w46436 & w40269;
	assign w40253 = w40270 & w40266;
	assign w14850 = ~w14853;
	assign w14951 = w14850 ^ w14851;
	assign w45305 = ~w14951;
	assign w43110 = w45305 ^ w45507;
	assign w50352 = w43165 ^ w43110;
	assign w46451 = w50352 ^ w417;
	assign w14136 = w46451 ^ w14140;
	assign w14123 = w14140 & w14136;
	assign w14053 = w46451 ^ w46449;
	assign w14134 = w14053 ^ w14142;
	assign w14143 = w46445 ^ w46451;
	assign w42978 = w43117 ^ w43110;
	assign w42977 = w42978 ^ w42979;
	assign w50360 = ~w42977;
	assign w42964 = w45305 ^ w32773;
	assign w50369 = w42963 ^ w42964;
	assign w42955 = w43076 ^ w45305;
	assign w50376 = w42954 ^ w42955;
	assign w42953 = w43112 ^ w43110;
	assign w46434 = w50369 ^ w434;
	assign w40200 = w46435 ^ w46434;
	assign w40265 = w40200 ^ w40267;
	assign w40268 = w40272 ^ w40200;
	assign w40274 = w46434 ^ w46432;
	assign w40259 = w40184 ^ w40274;
	assign w40271 = w46429 ^ w46434;
	assign w40250 = w40274 & w40259;
	assign w14133 = w46452 ^ w14134;
	assign w46443 = w50360 ^ w425;
	assign w10569 = w46443 ^ w46441;
	assign w10648 = w10569 ^ w10532;
	assign w10652 = w46443 ^ w10656;
	assign w10650 = w10569 ^ w10658;
	assign w10649 = w46444 ^ w10650;
	assign w46427 = w50376 ^ w441;
	assign w39596 = w46427 ^ w39600;
	assign w39603 = w46421 ^ w46427;
	assign w39583 = w39600 & w39596;
	assign w10639 = w10656 & w10652;
	assign w10659 = w46437 ^ w46443;
	assign w14132 = w14053 ^ w14016;
	assign w32786 = w32868 ^ w32885;
	assign w32781 = w32786 ^ w32882;
	assign w32860 = w32781 ^ w32784;
	assign w32847 = w32860 & w32892;
	assign w32825 = w32843 ^ w32847;
	assign w32803 = ~w32825;
	assign w32802 = w32803 ^ w32841;
	assign w32798 = w32802 ^ w44747;
	assign w32838 = w32860 & w32901;
	assign w32859 = w32781 ^ w32782;
	assign w32840 = w32859 & w32902;
	assign w43591 = w32839 ^ w32840;
	assign w32821 = w32845 ^ w43591;
	assign w32797 = w32821 ^ w32798;
	assign w50489 = w32796 ^ w32797;
	assign w43133 = w50484 ^ w50489;
	assign w42862 = ~w50489;
	assign w42937 = w42862 ^ w45293;
	assign w42909 = ~w43133;
	assign w42861 = w50495 ^ w42862;
	assign w32849 = w32859 & w32891;
	assign w32805 = w32848 ^ w32849;
	assign w32804 = w32849 ^ w32838;
	assign w32800 = ~w32804;
	assign w32822 = w32846 ^ w32821;
	assign w32826 = w32854 ^ w32822;
	assign w32831 = w32855 ^ w32826;
	assign w32795 = w32853 ^ w32826;
	assign w50491 = w44746 ^ w32831;
	assign w43118 = w50486 ^ w50491;
	assign w42906 = w50497 ^ w50491;
	assign w42890 = ~w43118;
	assign w42857 = w50491 ^ w50485;
	assign w32906 = w32831 ^ w32805;
	assign w50493 = ~w32906;
	assign w43104 = w45292 ^ w50493;
	assign w42929 = w32906 ^ w45291;
	assign w42901 = w45300 ^ w32906;
	assign w32801 = w32840 ^ w32798;
	assign w32905 = w32800 ^ w32801;
	assign w50492 = ~w32905;
	assign w43111 = w45291 ^ w50492;
	assign w42934 = w32905 ^ w50486;
	assign w42903 = w45299 ^ w32905;
	assign w32808 = w32812 ^ w43591;
	assign w32811 = w44747 ^ w32808;
	assign w32908 = w32810 ^ w32811;
	assign w50490 = w32794 ^ w32795;
	assign w43126 = w50485 ^ w50490;
	assign w42893 = ~w43126;
	assign w42855 = ~w50490;
	assign w42865 = w50496 ^ w42855;
	assign w42854 = w42855 ^ w50484;
	assign w32793 = w32849 ^ w32833;
	assign w50494 = w32822 ^ w32793;
	assign w43078 = w50487 ^ w50494;
	assign w43082 = w50494 ^ w50498;
	assign w42926 = w50494 ^ w45292;
	assign w42863 = ~w43082;
	assign w32807 = w32803 ^ w32808;
	assign w32907 = w32806 ^ w32807;
	assign w50488 = ~w32907;
	assign w43140 = w45293 ^ w50488;
	assign w42908 = w45301 ^ w32907;
	assign w42851 = w32907 ^ w45286;
	assign w45763 = ~w32908;
	assign w43141 = w45286 ^ w45763;
	assign w42910 = w43141 ^ w43082;
	assign w42859 = w45294 ^ w45763;
	assign w45899 = ~w43078;
	assign w42923 = w45899 ^ w45293;
	assign w42919 = w45899 ^ w50485;
	assign w42917 = w45899 ^ w50486;
	assign w14843 = w14888 ^ w14877;
	assign w14840 = ~w14843;
	assign w50476 = w14840 ^ w14841;
	assign w43107 = w50476 ^ w50480;
	assign w42990 = w43107 ^ w45507;
	assign w50353 = w42990 ^ w42991;
	assign w46450 = w50353 ^ w418;
	assign w14144 = w46450 ^ w46448;
	assign w14129 = w14054 ^ w14144;
	assign w14055 = w46450 ^ w14053;
	assign w14131 = w46446 ^ w14055;
	assign w14130 = w14060 ^ w14055;
	assign w14122 = w14137 & w14130;
	assign w14070 = w46451 ^ w46450;
	assign w14135 = w14070 ^ w14137;
	assign w14138 = w14142 ^ w14070;
	assign w14128 = w46447 ^ w14055;
	assign w14124 = w14143 & w14128;
	assign w14058 = w14124 ^ w14054;
	assign w14127 = w14134 & w14138;
	assign w14059 = w14127 ^ w14056;
	assign w14030 = w46449 ^ w46450;
	assign w14121 = w14142 & w14131;
	assign w14057 = w14121 ^ w14055;
	assign w14063 = w14059 ^ w14057;
	assign w14068 = w46445 ^ w14063;
	assign w42976 = w43116 ^ w43107;
	assign w50361 = w50467 ^ w42976;
	assign w46442 = w50361 ^ w426;
	assign w10571 = w46442 ^ w10569;
	assign w10586 = w46443 ^ w46442;
	assign w10657 = w46437 ^ w46442;
	assign w50377 = w50476 ^ w42953;
	assign w46426 = w50377 ^ w442;
	assign w39530 = w46427 ^ w46426;
	assign w39595 = w39530 ^ w39597;
	assign w39598 = w39602 ^ w39530;
	assign w39604 = w46426 ^ w46424;
	assign w39589 = w39514 ^ w39604;
	assign w39601 = w46421 ^ w46426;
	assign w39580 = w39604 & w39589;
	assign w42951 = w43109 ^ w43107;
	assign w50378 = w42951 ^ w42952;
	assign w46425 = w50378 ^ w443;
	assign w39513 = w46427 ^ w46425;
	assign w39515 = w46426 ^ w39513;
	assign w39591 = w46422 ^ w39515;
	assign w39588 = w46423 ^ w39515;
	assign w39590 = w39520 ^ w39515;
	assign w39594 = w39513 ^ w39602;
	assign w39593 = w46428 ^ w39594;
	assign w39490 = w46425 ^ w46426;
	assign w39592 = w39513 ^ w39476;
	assign w39587 = w39594 & w39598;
	assign w39519 = w39587 ^ w39516;
	assign w39586 = w39595 & w39593;
	assign w39537 = w39580 ^ w39586;
	assign w39584 = w39603 & w39588;
	assign w39518 = w39584 ^ w39514;
	assign w39582 = w39597 & w39590;
	assign w39581 = w39602 & w39591;
	assign w39517 = w39581 ^ w39515;
	assign w39523 = w39519 ^ w39517;
	assign w39528 = w46421 ^ w39523;
	assign w39578 = w39537 ^ w39528;
	assign w39489 = w39580 ^ w39581;
	assign w39536 = w39489 ^ w39490;
	assign w39535 = w39536 ^ w39518;
	assign w39577 = w39583 ^ w39535;
	assign w39579 = w39601 & w39592;
	assign w39574 = w39578 & w39577;
	assign w42846 = w50476 ^ w50472;
	assign w43159 = w42845 ^ w42846;
	assign w50370 = w43159 ^ w43109;
	assign w10644 = w46439 ^ w10571;
	assign w10640 = w10659 & w10644;
	assign w10574 = w10640 ^ w10570;
	assign w46433 = w50370 ^ w435;
	assign w40183 = w46435 ^ w46433;
	assign w40185 = w46434 ^ w40183;
	assign w40261 = w46430 ^ w40185;
	assign w40258 = w46431 ^ w40185;
	assign w40260 = w40190 ^ w40185;
	assign w40264 = w40183 ^ w40272;
	assign w40263 = w46436 ^ w40264;
	assign w40160 = w46433 ^ w46434;
	assign w40262 = w40183 ^ w40146;
	assign w40257 = w40264 & w40268;
	assign w40189 = w40257 ^ w40186;
	assign w40256 = w40265 & w40263;
	assign w40207 = w40250 ^ w40256;
	assign w40254 = w40273 & w40258;
	assign w40188 = w40254 ^ w40184;
	assign w40252 = w40267 & w40260;
	assign w40251 = w40272 & w40261;
	assign w40187 = w40251 ^ w40185;
	assign w40193 = w40189 ^ w40187;
	assign w40198 = w46429 ^ w40193;
	assign w40248 = w40207 ^ w40198;
	assign w40159 = w40250 ^ w40251;
	assign w40206 = w40159 ^ w40160;
	assign w40205 = w40206 ^ w40188;
	assign w40247 = w40253 ^ w40205;
	assign w40249 = w40271 & w40262;
	assign w40244 = w40248 & w40247;
	assign w10647 = w46438 ^ w10571;
	assign w14120 = w14144 & w14129;
	assign w14029 = w14120 ^ w14121;
	assign w14076 = w14029 ^ w14030;
	assign w14075 = w14076 ^ w14058;
	assign w14117 = w14123 ^ w14075;
	assign w10635 = w10657 & w10648;
	assign w10637 = w10658 & w10647;
	assign w10573 = w10637 ^ w10571;
	assign w10651 = w10586 ^ w10653;
	assign w10642 = w10651 & w10649;
	assign w10546 = w46441 ^ w46442;
	assign w10654 = w10658 ^ w10586;
	assign w45027 = w39579 ^ w39585;
	assign w39529 = w45027 ^ w39514;
	assign w39575 = w39537 ^ w39529;
	assign w39491 = w39523 ^ w45027;
	assign w39534 = w46423 ^ w39491;
	assign w39569 = w39574 ^ w39534;
	assign w45028 = w39579 ^ w39582;
	assign w39532 = w39580 ^ w45028;
	assign w39488 = w39583 ^ w39532;
	assign w39570 = w46427 ^ w39488;
	assign w39568 = w39569 & w39570;
	assign w39566 = w39574 ^ w39568;
	assign w39487 = w39568 ^ w39532;
	assign w39486 = w39568 ^ w39585;
	assign w39481 = w39486 ^ w39582;
	assign w39492 = w39518 ^ w45028;
	assign w39576 = w39492 ^ w39517;
	assign w39567 = w39568 ^ w39576;
	assign w39573 = w39574 ^ w39576;
	assign w39572 = w39575 & w39573;
	assign w39571 = w39572 ^ w39534;
	assign w39483 = w39572 ^ w39584;
	assign w39479 = w39483 ^ w39519;
	assign w39482 = w46421 ^ w39479;
	assign w39559 = w39481 ^ w39482;
	assign w39480 = w39572 ^ w39528;
	assign w39478 = w46423 ^ w39479;
	assign w39565 = w39576 & w39566;
	assign w39563 = w39565 ^ w39573;
	assign w39562 = w39571 & w39563;
	assign w39527 = w39562 ^ w39537;
	assign w39561 = w39527 ^ w39529;
	assign w39485 = w39562 ^ w39586;
	assign w39558 = w39527 ^ w39480;
	assign w39553 = w39567 & w46428;
	assign w39552 = w39558 & w39588;
	assign w39551 = w39561 & w39600;
	assign w39550 = w39571 & w39590;
	assign w39494 = w39550 ^ w39551;
	assign w39549 = w39559 & w39591;
	assign w39544 = w39567 & w39599;
	assign w39543 = w39558 & w39603;
	assign w39510 = w39552 ^ w39543;
	assign w39542 = w39561 & w39596;
	assign w39512 = w39550 ^ w39542;
	assign w39541 = w39571 & w39597;
	assign w39540 = w39559 & w39602;
	assign w45029 = w39551 ^ w39552;
	assign w45031 = w39565 ^ w39583;
	assign w39524 = w46427 ^ w45031;
	assign w39477 = w39524 ^ w39485;
	assign w39484 = w39514 ^ w39477;
	assign w39560 = w39481 ^ w39484;
	assign w39547 = w39560 & w39592;
	assign w39525 = w39543 ^ w39547;
	assign w39503 = ~w39525;
	assign w39556 = w39477 ^ w39478;
	assign w39548 = w39556 & w39589;
	assign w39509 = w39548 ^ w39551;
	assign w39506 = ~w39509;
	assign w39505 = w39548 ^ w39549;
	assign w39502 = w39503 ^ w39541;
	assign w39539 = w39556 & w39604;
	assign w39538 = w39560 & w39601;
	assign w39504 = w39549 ^ w39538;
	assign w39500 = ~w39504;
	assign w43608 = w39539 ^ w39540;
	assign w39508 = w39512 ^ w43608;
	assign w39507 = w39503 ^ w39508;
	assign w39607 = w39506 ^ w39507;
	assign w39533 = w39548 ^ w45029;
	assign w39499 = w39544 ^ w39533;
	assign w39496 = ~w39499;
	assign w39493 = w39549 ^ w39533;
	assign w39564 = w39524 ^ w39487;
	assign w39545 = w39564 & w39595;
	assign w39554 = w39564 & w39593;
	assign w39521 = w39545 ^ w43608;
	assign w39557 = w45031 ^ w39535;
	assign w39555 = w39557 & w39594;
	assign w39546 = w39557 & w39598;
	assign w39522 = w39546 ^ w39521;
	assign w39526 = w39554 ^ w39522;
	assign w39531 = w39555 ^ w39526;
	assign w50683 = w45029 ^ w39531;
	assign w39606 = w39531 ^ w39505;
	assign w39495 = w39553 ^ w39526;
	assign w50682 = w39494 ^ w39495;
	assign w50684 = w39522 ^ w39493;
	assign w45030 = w39553 ^ w39555;
	assign w39511 = w45030 ^ w39508;
	assign w39608 = w39510 ^ w39511;
	assign w39498 = w39502 ^ w45030;
	assign w39501 = w39540 ^ w39498;
	assign w39605 = w39500 ^ w39501;
	assign w39497 = w39521 ^ w39498;
	assign w50681 = w39496 ^ w39497;
	assign w45055 = w40249 ^ w40252;
	assign w40162 = w40188 ^ w45055;
	assign w40246 = w40162 ^ w40187;
	assign w40243 = w40244 ^ w40246;
	assign w40202 = w40250 ^ w45055;
	assign w40158 = w40253 ^ w40202;
	assign w40240 = w46435 ^ w40158;
	assign w45058 = w40249 ^ w40255;
	assign w40161 = w40193 ^ w45058;
	assign w40204 = w46431 ^ w40161;
	assign w40239 = w40244 ^ w40204;
	assign w40238 = w40239 & w40240;
	assign w40236 = w40244 ^ w40238;
	assign w40157 = w40238 ^ w40202;
	assign w40156 = w40238 ^ w40255;
	assign w40151 = w40156 ^ w40252;
	assign w40235 = w40246 & w40236;
	assign w40233 = w40235 ^ w40243;
	assign w45057 = w40235 ^ w40253;
	assign w40227 = w45057 ^ w40205;
	assign w40216 = w40227 & w40268;
	assign w40225 = w40227 & w40264;
	assign w40194 = w46435 ^ w45057;
	assign w40234 = w40194 ^ w40157;
	assign w40224 = w40234 & w40263;
	assign w40215 = w40234 & w40265;
	assign w40237 = w40238 ^ w40246;
	assign w40223 = w40237 & w46436;
	assign w40214 = w40237 & w40269;
	assign w40199 = w45058 ^ w40184;
	assign w40245 = w40207 ^ w40199;
	assign w40242 = w40245 & w40243;
	assign w40241 = w40242 ^ w40204;
	assign w40153 = w40242 ^ w40254;
	assign w40149 = w40153 ^ w40189;
	assign w40152 = w46429 ^ w40149;
	assign w40229 = w40151 ^ w40152;
	assign w40150 = w40242 ^ w40198;
	assign w40148 = w46431 ^ w40149;
	assign w40232 = w40241 & w40233;
	assign w40197 = w40232 ^ w40207;
	assign w40231 = w40197 ^ w40199;
	assign w40155 = w40232 ^ w40256;
	assign w40147 = w40194 ^ w40155;
	assign w40154 = w40184 ^ w40147;
	assign w40230 = w40151 ^ w40154;
	assign w40228 = w40197 ^ w40150;
	assign w40226 = w40147 ^ w40148;
	assign w40222 = w40228 & w40258;
	assign w40221 = w40231 & w40270;
	assign w40220 = w40241 & w40260;
	assign w40164 = w40220 ^ w40221;
	assign w40219 = w40229 & w40261;
	assign w40218 = w40226 & w40259;
	assign w40179 = w40218 ^ w40221;
	assign w40176 = ~w40179;
	assign w40175 = w40218 ^ w40219;
	assign w40217 = w40230 & w40262;
	assign w40213 = w40228 & w40273;
	assign w40195 = w40213 ^ w40217;
	assign w40180 = w40222 ^ w40213;
	assign w40173 = ~w40195;
	assign w40212 = w40231 & w40266;
	assign w40182 = w40220 ^ w40212;
	assign w40211 = w40241 & w40267;
	assign w40172 = w40173 ^ w40211;
	assign w40210 = w40229 & w40272;
	assign w40209 = w40226 & w40274;
	assign w40208 = w40230 & w40271;
	assign w40174 = w40219 ^ w40208;
	assign w40170 = ~w40174;
	assign w45056 = w40209 ^ w40210;
	assign w40191 = w40215 ^ w45056;
	assign w40192 = w40216 ^ w40191;
	assign w40196 = w40224 ^ w40192;
	assign w40165 = w40223 ^ w40196;
	assign w50697 = w40164 ^ w40165;
	assign w40201 = w40225 ^ w40196;
	assign w40276 = w40201 ^ w40175;
	assign w40178 = w40182 ^ w45056;
	assign w40177 = w40173 ^ w40178;
	assign w40277 = w40176 ^ w40177;
	assign w45059 = w40221 ^ w40222;
	assign w50698 = w45059 ^ w40201;
	assign w40203 = w40218 ^ w45059;
	assign w40169 = w40214 ^ w40203;
	assign w40166 = ~w40169;
	assign w40163 = w40219 ^ w40203;
	assign w50699 = w40192 ^ w40163;
	assign w45060 = w40223 ^ w40225;
	assign w40181 = w45060 ^ w40178;
	assign w40278 = w40180 ^ w40181;
	assign w40168 = w40172 ^ w45060;
	assign w40171 = w40210 ^ w40168;
	assign w40275 = w40170 ^ w40171;
	assign w40167 = w40191 ^ w40168;
	assign w50696 = w40166 ^ w40167;
	assign w14141 = w46445 ^ w46450;
	assign w14119 = w14141 & w14132;
	assign w43958 = w14119 ^ w14122;
	assign w14032 = w14058 ^ w43958;
	assign w14116 = w14032 ^ w14057;
	assign w14072 = w14120 ^ w43958;
	assign w14028 = w14123 ^ w14072;
	assign w14110 = w46451 ^ w14028;
	assign w43961 = w14119 ^ w14125;
	assign w14031 = w14063 ^ w43961;
	assign w14074 = w46447 ^ w14031;
	assign w14069 = w43961 ^ w14054;
	assign w10643 = w10650 & w10654;
	assign w10575 = w10643 ^ w10572;
	assign w10579 = w10575 ^ w10573;
	assign w10584 = w46437 ^ w10579;
	assign w43814 = w10635 ^ w10641;
	assign w10547 = w10579 ^ w43814;
	assign w10590 = w46439 ^ w10547;
	assign w10585 = w43814 ^ w10570;
	assign w10646 = w10576 ^ w10571;
	assign w10638 = w10653 & w10646;
	assign w43815 = w10635 ^ w10638;
	assign w10548 = w10574 ^ w43815;
	assign w10632 = w10548 ^ w10573;
	assign w45818 = ~w39606;
	assign w45819 = ~w39607;
	assign w45820 = ~w39608;
	assign w45825 = ~w39605;
	assign w45834 = ~w40276;
	assign w45835 = ~w40277;
	assign w45836 = ~w40278;
	assign w45841 = ~w40275;
	assign w14126 = w14135 & w14133;
	assign w14077 = w14120 ^ w14126;
	assign w14118 = w14077 ^ w14068;
	assign w14114 = w14118 & w14117;
	assign w14113 = w14114 ^ w14116;
	assign w14109 = w14114 ^ w14074;
	assign w14108 = w14109 & w14110;
	assign w14107 = w14108 ^ w14116;
	assign w14026 = w14108 ^ w14125;
	assign w14021 = w14026 ^ w14122;
	assign w14106 = w14114 ^ w14108;
	assign w14105 = w14116 & w14106;
	assign w14103 = w14105 ^ w14113;
	assign w43960 = w14105 ^ w14123;
	assign w14097 = w43960 ^ w14075;
	assign w14095 = w14097 & w14134;
	assign w14086 = w14097 & w14138;
	assign w14064 = w46451 ^ w43960;
	assign w14093 = w14107 & w46452;
	assign w43963 = w14093 ^ w14095;
	assign w14084 = w14107 & w14139;
	assign w14027 = w14108 ^ w14072;
	assign w14104 = w14064 ^ w14027;
	assign w14094 = w14104 & w14133;
	assign w14115 = w14077 ^ w14069;
	assign w14112 = w14115 & w14113;
	assign w14023 = w14112 ^ w14124;
	assign w14111 = w14112 ^ w14074;
	assign w14019 = w14023 ^ w14059;
	assign w14102 = w14111 & w14103;
	assign w14025 = w14102 ^ w14126;
	assign w14017 = w14064 ^ w14025;
	assign w14024 = w14054 ^ w14017;
	assign w14090 = w14111 & w14130;
	assign w14081 = w14111 & w14137;
	assign w14100 = w14021 ^ w14024;
	assign w14078 = w14100 & w14141;
	assign w14087 = w14100 & w14132;
	assign w14022 = w46445 ^ w14019;
	assign w14099 = w14021 ^ w14022;
	assign w14080 = w14099 & w14142;
	assign w14089 = w14099 & w14131;
	assign w14044 = w14089 ^ w14078;
	assign w14040 = ~w14044;
	assign w14067 = w14102 ^ w14077;
	assign w14101 = w14067 ^ w14069;
	assign w14091 = w14101 & w14140;
	assign w14034 = w14090 ^ w14091;
	assign w14020 = w14112 ^ w14068;
	assign w14098 = w14067 ^ w14020;
	assign w14092 = w14098 & w14128;
	assign w14083 = w14098 & w14143;
	assign w43962 = w14091 ^ w14092;
	assign w14050 = w14092 ^ w14083;
	assign w14065 = w14083 ^ w14087;
	assign w14043 = ~w14065;
	assign w14042 = w14043 ^ w14081;
	assign w14038 = w14042 ^ w43963;
	assign w14041 = w14080 ^ w14038;
	assign w14145 = w14040 ^ w14041;
	assign w14018 = w46447 ^ w14019;
	assign w14096 = w14017 ^ w14018;
	assign w14079 = w14096 & w14144;
	assign w43959 = w14079 ^ w14080;
	assign w14088 = w14096 & w14129;
	assign w14049 = w14088 ^ w14091;
	assign w14073 = w14088 ^ w43962;
	assign w14039 = w14084 ^ w14073;
	assign w14036 = ~w14039;
	assign w14033 = w14089 ^ w14073;
	assign w14046 = ~w14049;
	assign w14045 = w14088 ^ w14089;
	assign w45278 = ~w14145;
	assign w14085 = w14104 & w14135;
	assign w14061 = w14085 ^ w43959;
	assign w14062 = w14086 ^ w14061;
	assign w14037 = w14061 ^ w14038;
	assign w50651 = w14062 ^ w14033;
	assign w14066 = w14094 ^ w14062;
	assign w14071 = w14095 ^ w14066;
	assign w14035 = w14093 ^ w14066;
	assign w14146 = w14071 ^ w14045;
	assign w50649 = w14034 ^ w14035;
	assign w50648 = w14036 ^ w14037;
	assign w50650 = w43962 ^ w14071;
	assign w45279 = ~w14146;
	assign w14082 = w14101 & w14136;
	assign w14052 = w14090 ^ w14082;
	assign w14048 = w14052 ^ w43959;
	assign w14051 = w43963 ^ w14048;
	assign w14047 = w14043 ^ w14048;
	assign w14148 = w14050 ^ w14051;
	assign w14147 = w14046 ^ w14047;
	assign w45280 = ~w14147;
	assign w45281 = ~w14148;
	assign w10660 = w46442 ^ w46440;
	assign w10645 = w10570 ^ w10660;
	assign w10636 = w10660 & w10645;
	assign w10593 = w10636 ^ w10642;
	assign w10631 = w10593 ^ w10585;
	assign w10545 = w10636 ^ w10637;
	assign w10592 = w10545 ^ w10546;
	assign w10591 = w10592 ^ w10574;
	assign w10633 = w10639 ^ w10591;
	assign w10588 = w10636 ^ w43815;
	assign w10544 = w10639 ^ w10588;
	assign w10626 = w46443 ^ w10544;
	assign w10634 = w10593 ^ w10584;
	assign w10630 = w10634 & w10633;
	assign w10625 = w10630 ^ w10590;
	assign w10629 = w10630 ^ w10632;
	assign w10628 = w10631 & w10629;
	assign w10627 = w10628 ^ w10590;
	assign w10606 = w10627 & w10646;
	assign w10539 = w10628 ^ w10640;
	assign w10535 = w10539 ^ w10575;
	assign w10534 = w46439 ^ w10535;
	assign w10624 = w10625 & w10626;
	assign w10623 = w10624 ^ w10632;
	assign w10542 = w10624 ^ w10641;
	assign w10622 = w10630 ^ w10624;
	assign w10621 = w10632 & w10622;
	assign w10619 = w10621 ^ w10629;
	assign w10618 = w10627 & w10619;
	assign w10541 = w10618 ^ w10642;
	assign w10537 = w10542 ^ w10638;
	assign w10600 = w10623 & w10655;
	assign w10609 = w10623 & w46444;
	assign w43818 = w10621 ^ w10639;
	assign w10580 = w46443 ^ w43818;
	assign w10597 = w10627 & w10653;
	assign w10583 = w10618 ^ w10593;
	assign w10613 = w43818 ^ w10591;
	assign w10611 = w10613 & w10650;
	assign w10533 = w10580 ^ w10541;
	assign w10612 = w10533 ^ w10534;
	assign w10595 = w10612 & w10660;
	assign w10604 = w10612 & w10645;
	assign w10536 = w10628 ^ w10584;
	assign w10543 = w10624 ^ w10588;
	assign w10620 = w10580 ^ w10543;
	assign w10610 = w10620 & w10649;
	assign w10601 = w10620 & w10651;
	assign w10602 = w10613 & w10654;
	assign w10538 = w46437 ^ w10535;
	assign w10615 = w10537 ^ w10538;
	assign w10605 = w10615 & w10647;
	assign w10614 = w10583 ^ w10536;
	assign w10599 = w10614 & w10659;
	assign w10608 = w10614 & w10644;
	assign w10566 = w10608 ^ w10599;
	assign w10596 = w10615 & w10658;
	assign w43525 = w10595 ^ w10596;
	assign w10577 = w10601 ^ w43525;
	assign w43817 = w10609 ^ w10611;
	assign w10540 = w10570 ^ w10533;
	assign w10616 = w10537 ^ w10540;
	assign w10603 = w10616 & w10648;
	assign w10594 = w10616 & w10657;
	assign w10560 = w10605 ^ w10594;
	assign w10556 = ~w10560;
	assign w10581 = w10599 ^ w10603;
	assign w10559 = ~w10581;
	assign w10558 = w10559 ^ w10597;
	assign w10554 = w10558 ^ w43817;
	assign w10557 = w10596 ^ w10554;
	assign w10661 = w10556 ^ w10557;
	assign w10553 = w10577 ^ w10554;
	assign w45215 = ~w10661;
	assign w10617 = w10583 ^ w10585;
	assign w10607 = w10617 & w10656;
	assign w10550 = w10606 ^ w10607;
	assign w10598 = w10617 & w10652;
	assign w10568 = w10606 ^ w10598;
	assign w10565 = w10604 ^ w10607;
	assign w10562 = ~w10565;
	assign w10564 = w10568 ^ w43525;
	assign w10563 = w10559 ^ w10564;
	assign w10567 = w43817 ^ w10564;
	assign w10664 = w10566 ^ w10567;
	assign w10663 = w10562 ^ w10563;
	assign w45213 = ~w10664;
	assign w45217 = ~w10663;
	assign w43816 = w10607 ^ w10608;
	assign w10589 = w10604 ^ w43816;
	assign w10549 = w10605 ^ w10589;
	assign w10555 = w10600 ^ w10589;
	assign w10552 = ~w10555;
	assign w50709 = w10552 ^ w10553;
	assign w10561 = w10604 ^ w10605;
	assign w10578 = w10602 ^ w10577;
	assign w50712 = w10578 ^ w10549;
	assign w10582 = w10610 ^ w10578;
	assign w10587 = w10611 ^ w10582;
	assign w10662 = w10587 ^ w10561;
	assign w10551 = w10609 ^ w10582;
	assign w50710 = w10550 ^ w10551;
	assign w50711 = w43816 ^ w10587;
	assign w9792 = w45215 ^ w50711;
	assign w45216 = ~w10662;
	assign w9577 = w50710 ^ w50709;
	assign w45970 = ~w43423;
	assign w43342 = w45970 ^ w50259;
	assign w50146 = w43341 ^ w43342;
	assign w46584 = w50146 ^ w1337;
	assign w29332 = w46584 ^ w46582;
	assign w29291 = w29332 ^ w46583;
	assign w29415 = w46588 ^ w29291;
	assign w29292 = w29332 ^ w29330;
	assign w43255 = w45970 ^ w45325;
	assign w50125 = w43255 ^ w43256;
	assign w46605 = w50125 ^ w1316;
	assign w15079 = w46605 ^ w46610;
	assign w43218 = w45970 ^ w50261;
	assign w43491 = w43218 ^ w43219;
	assign w50145 = w43491 ^ w43488;
	assign w29401 = w46588 & w29415;
	assign w29418 = w46584 ^ w46581;
	assign w46585 = w50145 ^ w1336;
	assign w29306 = w46585 ^ w46586;
	assign w14992 = w46607 ^ w46605;
	assign w14954 = w14994 ^ w14992;
	assign w15075 = w14992 ^ w14998;
	assign w15073 = w15008 ^ w15075;
	assign w15060 = w15075 & w15068;
	assign w15067 = w14992 ^ w15082;
	assign w15058 = w15082 & w15067;
	assign w15081 = w46605 ^ w46611;
	assign w15062 = w15081 & w15066;
	assign w14996 = w15062 ^ w14992;
	assign w29414 = w29418 ^ w29346;
	assign w15080 = w46608 ^ w46605;
	assign w15076 = w15080 ^ w15008;
	assign w15059 = w15080 & w15069;
	assign w14995 = w15059 ^ w14993;
	assign w15072 = w14991 ^ w15080;
	assign w15065 = w15072 & w15076;
	assign w14997 = w15065 ^ w14994;
	assign w15071 = w46612 ^ w15072;
	assign w15064 = w15073 & w15071;
	assign w15001 = w14997 ^ w14995;
	assign w14967 = w15058 ^ w15059;
	assign w15014 = w14967 ^ w14968;
	assign w15013 = w15014 ^ w14996;
	assign w15055 = w15061 ^ w15013;
	assign w15015 = w15058 ^ w15064;
	assign w15070 = w14991 ^ w14954;
	assign w15057 = w15079 & w15070;
	assign w43997 = w15057 ^ w15060;
	assign w14970 = w14996 ^ w43997;
	assign w15054 = w14970 ^ w14995;
	assign w44000 = w15057 ^ w15063;
	assign w15010 = w15058 ^ w43997;
	assign w14966 = w15061 ^ w15010;
	assign w15007 = w44000 ^ w14992;
	assign w15053 = w15015 ^ w15007;
	assign w15048 = w46611 ^ w14966;
	assign w14969 = w15001 ^ w44000;
	assign w15012 = w46607 ^ w14969;
	assign w29420 = w46586 ^ w46584;
	assign w29405 = w29330 ^ w29420;
	assign w29396 = w29420 & w29405;
	assign w29329 = w46587 ^ w46585;
	assign w29331 = w46586 ^ w29329;
	assign w29407 = w46582 ^ w29331;
	assign w29408 = w29329 ^ w29292;
	assign w29404 = w46583 ^ w29331;
	assign w29400 = w29419 & w29404;
	assign w29334 = w29400 ^ w29330;
	assign w29410 = w29329 ^ w29418;
	assign w29403 = w29410 & w29414;
	assign w29335 = w29403 ^ w29332;
	assign w29409 = w46588 ^ w29410;
	assign w29402 = w29411 & w29409;
	assign w29395 = w29417 & w29408;
	assign w44598 = w29395 ^ w29401;
	assign w29345 = w44598 ^ w29330;
	assign w29353 = w29396 ^ w29402;
	assign w29391 = w29353 ^ w29345;
	assign w29406 = w29336 ^ w29331;
	assign w29398 = w29413 & w29406;
	assign w44599 = w29395 ^ w29398;
	assign w29348 = w29396 ^ w44599;
	assign w29304 = w29399 ^ w29348;
	assign w29308 = w29334 ^ w44599;
	assign w29386 = w46587 ^ w29304;
	assign w29397 = w29418 & w29407;
	assign w29305 = w29396 ^ w29397;
	assign w29333 = w29397 ^ w29331;
	assign w29392 = w29308 ^ w29333;
	assign w29352 = w29305 ^ w29306;
	assign w29339 = w29335 ^ w29333;
	assign w29344 = w46581 ^ w29339;
	assign w29394 = w29353 ^ w29344;
	assign w29307 = w29339 ^ w44598;
	assign w29350 = w46583 ^ w29307;
	assign w29351 = w29352 ^ w29334;
	assign w29393 = w29399 ^ w29351;
	assign w29390 = w29394 & w29393;
	assign w29389 = w29390 ^ w29392;
	assign w29385 = w29390 ^ w29350;
	assign w29388 = w29391 & w29389;
	assign w29299 = w29388 ^ w29400;
	assign w29295 = w29299 ^ w29335;
	assign w29294 = w46583 ^ w29295;
	assign w29296 = w29388 ^ w29344;
	assign w29298 = w46581 ^ w29295;
	assign w29384 = w29385 & w29386;
	assign w29382 = w29390 ^ w29384;
	assign w29303 = w29384 ^ w29348;
	assign w29383 = w29384 ^ w29392;
	assign w29369 = w29383 & w46588;
	assign w29360 = w29383 & w29415;
	assign w29302 = w29384 ^ w29401;
	assign w29297 = w29302 ^ w29398;
	assign w29375 = w29297 ^ w29298;
	assign w29356 = w29375 & w29418;
	assign w29365 = w29375 & w29407;
	assign w29387 = w29388 ^ w29350;
	assign w29357 = w29387 & w29413;
	assign w29366 = w29387 & w29406;
	assign w29381 = w29392 & w29382;
	assign w29379 = w29381 ^ w29389;
	assign w29378 = w29387 & w29379;
	assign w44602 = w29381 ^ w29399;
	assign w29340 = w46587 ^ w44602;
	assign w29380 = w29340 ^ w29303;
	assign w29370 = w29380 & w29409;
	assign w29361 = w29380 & w29411;
	assign w29373 = w44602 ^ w29351;
	assign w29371 = w29373 & w29410;
	assign w29362 = w29373 & w29414;
	assign w44601 = w29369 ^ w29371;
	assign w29343 = w29378 ^ w29353;
	assign w29374 = w29343 ^ w29296;
	assign w29359 = w29374 & w29419;
	assign w29368 = w29374 & w29404;
	assign w29377 = w29343 ^ w29345;
	assign w29358 = w29377 & w29412;
	assign w29326 = w29368 ^ w29359;
	assign w29367 = w29377 & w29416;
	assign w29310 = w29366 ^ w29367;
	assign w29328 = w29366 ^ w29358;
	assign w44600 = w29367 ^ w29368;
	assign w29301 = w29378 ^ w29402;
	assign w29293 = w29340 ^ w29301;
	assign w29372 = w29293 ^ w29294;
	assign w29300 = w29330 ^ w29293;
	assign w29364 = w29372 & w29405;
	assign w29325 = w29364 ^ w29367;
	assign w29321 = w29364 ^ w29365;
	assign w29322 = ~w29325;
	assign w29349 = w29364 ^ w44600;
	assign w29309 = w29365 ^ w29349;
	assign w29315 = w29360 ^ w29349;
	assign w29312 = ~w29315;
	assign w29355 = w29372 & w29420;
	assign w43581 = w29355 ^ w29356;
	assign w29337 = w29361 ^ w43581;
	assign w29338 = w29362 ^ w29337;
	assign w29342 = w29370 ^ w29338;
	assign w29311 = w29369 ^ w29342;
	assign w50463 = w29310 ^ w29311;
	assign w43134 = w50459 ^ w50463;
	assign w50330 = w43149 ^ w43134;
	assign w46473 = w50330 ^ w459;
	assign w43014 = w43015 ^ w50463;
	assign w50338 = w43013 ^ w43014;
	assign w42999 = w43135 ^ w43134;
	assign w42997 = ~w42999;
	assign w42830 = w50463 ^ w50453;
	assign w29347 = w29371 ^ w29342;
	assign w29422 = w29347 ^ w29321;
	assign w42912 = w29422 ^ w50456;
	assign w43006 = w43130 ^ w29422;
	assign w50341 = w43006 ^ w43007;
	assign w29324 = w29328 ^ w43581;
	assign w50465 = ~w29422;
	assign w43124 = w45288 ^ w50465;
	assign w43022 = w43132 ^ w43124;
	assign w50333 = w45584 ^ w43022;
	assign w46470 = w50333 ^ w462;
	assign w42993 = w43124 ^ w43080;
	assign w50350 = w50461 ^ w42993;
	assign w42931 = w43124 ^ w45583;
	assign w46453 = w50350 ^ w479;
	assign w29327 = w44601 ^ w29324;
	assign w29424 = w29326 ^ w29327;
	assign w46465 = w50338 ^ w467;
	assign w50466 = w29338 ^ w29309;
	assign w43079 = w50461 ^ w50466;
	assign w43087 = w50450 ^ w50466;
	assign w43072 = w43120 ^ w43087;
	assign w43021 = w43130 ^ w43079;
	assign w50334 = w50450 ^ w43021;
	assign w42983 = ~w43087;
	assign w43004 = w45964 ^ w50466;
	assign w50342 = w43004 ^ w43005;
	assign w43003 = w43120 ^ w43079;
	assign w50343 = w45578 ^ w43003;
	assign w42982 = w42983 ^ w50452;
	assign w42829 = w43087 ^ w50448;
	assign w43166 = w42829 ^ w42830;
	assign w46461 = w50342 ^ w471;
	assign w46460 = w50343 ^ w472;
	assign w46469 = w50334 ^ w463;
	assign w45667 = ~w29424;
	assign w43143 = w45578 ^ w45667;
	assign w50319 = w45667 ^ w43072;
	assign w43020 = w43143 ^ w43081;
	assign w50335 = w45221 ^ w43020;
	assign w43011 = w43143 ^ w43121;
	assign w42895 = w43143 ^ w43080;
	assign w50327 = w45289 ^ w42895;
	assign w46476 = w50327 ^ w456;
	assign w42872 = w43079 ^ w45667;
	assign w43148 = w42872 ^ w42873;
	assign w50344 = w43148 ^ w43121;
	assign w46484 = w50319 ^ w448;
	assign w46459 = w50344 ^ w473;
	assign w23523 = w46453 ^ w46459;
	assign w10710 = w46476 ^ w46470;
	assign w46468 = w50335 ^ w464;
	assign w29376 = w29297 ^ w29300;
	assign w29363 = w29376 & w29408;
	assign w29354 = w29376 & w29417;
	assign w29320 = w29365 ^ w29354;
	assign w29316 = ~w29320;
	assign w29341 = w29359 ^ w29363;
	assign w29319 = ~w29341;
	assign w29323 = w29319 ^ w29324;
	assign w29423 = w29322 ^ w29323;
	assign w45666 = ~w29423;
	assign w43142 = w45585 ^ w45666;
	assign w50328 = w43150 ^ w43142;
	assign w46475 = w50328 ^ w457;
	assign w10793 = w46469 ^ w46475;
	assign w10703 = w46475 ^ w46473;
	assign w43018 = w43142 ^ w43120;
	assign w43017 = w43018 ^ w43019;
	assign w50336 = ~w43017;
	assign w43012 = w42983 ^ w45666;
	assign w43010 = w43011 ^ w43012;
	assign w50320 = ~w43010;
	assign w43001 = w45666 ^ w14415;
	assign w50345 = w43000 ^ w43001;
	assign w46458 = w50345 ^ w474;
	assign w42995 = w43142 ^ w43119;
	assign w46483 = w50320 ^ w449;
	assign w23450 = w46459 ^ w46458;
	assign w46467 = w50336 ^ w465;
	assign w14277 = w46461 ^ w46467;
	assign w14187 = w46467 ^ w46465;
	assign w23521 = w46453 ^ w46458;
	assign w46462 = w50341 ^ w470;
	assign w14194 = w46468 ^ w46462;
	assign w50464 = w44600 ^ w29347;
	assign w43131 = w50460 ^ w50464;
	assign w50323 = w43166 ^ w43131;
	assign w46480 = w50323 ^ w452;
	assign w43024 = w43026 ^ w43131;
	assign w50331 = w43024 ^ w43025;
	assign w42996 = w43132 ^ w43131;
	assign w50348 = w45287 ^ w42996;
	assign w42949 = w50464 ^ w10929;
	assign w46472 = w50331 ^ w460;
	assign w42866 = w43081 ^ w50464;
	assign w43151 = w42866 ^ w42867;
	assign w50339 = w43151 ^ w43135;
	assign w46455 = w50348 ^ w477;
	assign w23434 = w46455 ^ w46453;
	assign w10792 = w46472 ^ w46469;
	assign w10784 = w10703 ^ w10792;
	assign w10783 = w46476 ^ w10784;
	assign w46464 = w50339 ^ w468;
	assign w14276 = w46464 ^ w46461;
	assign w14268 = w14187 ^ w14276;
	assign w14190 = w46464 ^ w46462;
	assign w14267 = w46468 ^ w14268;
	assign w10706 = w46472 ^ w46470;
	assign w29318 = w29319 ^ w29357;
	assign w29314 = w29318 ^ w44601;
	assign w29317 = w29356 ^ w29314;
	assign w29421 = w29316 ^ w29317;
	assign w29313 = w29337 ^ w29314;
	assign w50462 = w29312 ^ w29313;
	assign w43122 = w50447 ^ w50462;
	assign w42984 = ~w43122;
	assign w43053 = w42984 ^ w45220;
	assign w50329 = w43053 ^ w43054;
	assign w43016 = w43122 ^ w43121;
	assign w50337 = w50451 ^ w43016;
	assign w46466 = w50337 ^ w466;
	assign w14204 = w46467 ^ w46466;
	assign w14164 = w46465 ^ w46466;
	assign w14272 = w14276 ^ w14204;
	assign w14189 = w46466 ^ w14187;
	assign w14265 = w46462 ^ w14189;
	assign w14255 = w14276 & w14265;
	assign w14261 = w14268 & w14272;
	assign w14278 = w46466 ^ w46464;
	assign w50321 = w50462 ^ w42995;
	assign w42981 = w43134 ^ w42984;
	assign w50322 = w42981 ^ w42982;
	assign w14264 = w14194 ^ w14189;
	assign w14275 = w46461 ^ w46466;
	assign w14191 = w14255 ^ w14189;
	assign w46482 = w50321 ^ w450;
	assign w25996 = w46483 ^ w46482;
	assign w26070 = w46482 ^ w46480;
	assign w14193 = w14261 ^ w14190;
	assign w14197 = w14193 ^ w14191;
	assign w14202 = w46461 ^ w14197;
	assign w46474 = w50329 ^ w458;
	assign w10720 = w46475 ^ w46474;
	assign w10680 = w46473 ^ w46474;
	assign w10791 = w46469 ^ w46474;
	assign w10794 = w46474 ^ w46472;
	assign w10705 = w46474 ^ w10703;
	assign w10780 = w10710 ^ w10705;
	assign w10788 = w10792 ^ w10720;
	assign w10777 = w10784 & w10788;
	assign w10709 = w10777 ^ w10706;
	assign w45673 = ~w29421;
	assign w43127 = w45287 ^ w45673;
	assign w43023 = w43135 ^ w43127;
	assign w50332 = w45583 ^ w43023;
	assign w43008 = w43132 ^ w45673;
	assign w50340 = w43008 ^ w43009;
	assign w46463 = w50340 ^ w469;
	assign w42994 = w43130 ^ w43127;
	assign w50349 = w45288 ^ w42994;
	assign w46454 = w50349 ^ w478;
	assign w23440 = w46460 ^ w46454;
	assign w23520 = w46455 ^ w23440;
	assign w42950 = w43127 ^ w50449;
	assign w42948 = ~w42950;
	assign w50324 = w42948 ^ w42949;
	assign w42932 = w45673 ^ w10930;
	assign w42930 = w42931 ^ w42932;
	assign w50325 = ~w42930;
	assign w46478 = w50325 ^ w454;
	assign w46471 = w50332 ^ w461;
	assign w10665 = w10706 ^ w46471;
	assign w10790 = w46471 ^ w10710;
	assign w14188 = w46463 ^ w46461;
	assign w14150 = w14190 ^ w14188;
	assign w14262 = w46463 ^ w14189;
	assign w14258 = w14277 & w14262;
	assign w14274 = w46463 ^ w14194;
	assign w14270 = w46467 ^ w14274;
	assign w14257 = w14274 & w14270;
	assign w25982 = w46480 ^ w46478;
	assign w25986 = w46484 ^ w46478;
	assign w23517 = w23434 ^ w23440;
	assign w23515 = w23450 ^ w23517;
	assign w10704 = w46471 ^ w46469;
	assign w10787 = w10704 ^ w10710;
	assign w10785 = w10720 ^ w10787;
	assign w10776 = w10785 & w10783;
	assign w10666 = w10706 ^ w10704;
	assign w10782 = w10703 ^ w10666;
	assign w10769 = w10791 & w10782;
	assign w10772 = w10787 & w10780;
	assign w14271 = w14188 ^ w14194;
	assign w14256 = w14271 & w14264;
	assign w14266 = w14187 ^ w14150;
	assign w14253 = w14275 & w14266;
	assign w43965 = w14253 ^ w14256;
	assign w10789 = w46476 ^ w10665;
	assign w10775 = w46476 & w10789;
	assign w43819 = w10769 ^ w10775;
	assign w10719 = w43819 ^ w10704;
	assign w14192 = w14258 ^ w14188;
	assign w14166 = w14192 ^ w43965;
	assign w14250 = w14166 ^ w14191;
	assign w10778 = w46471 ^ w10705;
	assign w10774 = w10793 & w10778;
	assign w10708 = w10774 ^ w10704;
	assign w10779 = w10704 ^ w10794;
	assign w10770 = w10794 & w10779;
	assign w10727 = w10770 ^ w10776;
	assign w10765 = w10727 ^ w10719;
	assign w46479 = w50324 ^ w453;
	assign w14149 = w14190 ^ w46463;
	assign w14273 = w46468 ^ w14149;
	assign w14259 = w46468 & w14273;
	assign w43964 = w14253 ^ w14259;
	assign w14165 = w14197 ^ w43964;
	assign w14203 = w43964 ^ w14188;
	assign w26066 = w46479 ^ w25986;
	assign w26062 = w46483 ^ w26066;
	assign w26049 = w26066 & w26062;
	assign w10786 = w46475 ^ w10790;
	assign w10773 = w10790 & w10786;
	assign w43820 = w10769 ^ w10772;
	assign w10682 = w10708 ^ w43820;
	assign w10722 = w10770 ^ w43820;
	assign w10678 = w10773 ^ w10722;
	assign w10760 = w46475 ^ w10678;
	assign w14263 = w14188 ^ w14278;
	assign w14254 = w14278 & w14263;
	assign w14163 = w14254 ^ w14255;
	assign w14210 = w14163 ^ w14164;
	assign w14209 = w14210 ^ w14192;
	assign w14251 = w14257 ^ w14209;
	assign w14206 = w14254 ^ w43965;
	assign w14162 = w14257 ^ w14206;
	assign w14244 = w46467 ^ w14162;
	assign w25941 = w25982 ^ w46479;
	assign w26065 = w46484 ^ w25941;
	assign w26051 = w46484 & w26065;
	assign w14269 = w14204 ^ w14271;
	assign w14260 = w14269 & w14267;
	assign w14211 = w14254 ^ w14260;
	assign w14252 = w14211 ^ w14202;
	assign w14248 = w14252 & w14251;
	assign w14247 = w14248 ^ w14250;
	assign w14249 = w14211 ^ w14203;
	assign w14246 = w14249 & w14247;
	assign w14154 = w14246 ^ w14202;
	assign w14157 = w14246 ^ w14258;
	assign w14153 = w14157 ^ w14193;
	assign w14152 = w46463 ^ w14153;
	assign w14156 = w46461 ^ w14153;
	assign w10781 = w46470 ^ w10705;
	assign w10771 = w10792 & w10781;
	assign w10679 = w10770 ^ w10771;
	assign w10726 = w10679 ^ w10680;
	assign w10725 = w10726 ^ w10708;
	assign w10767 = w10773 ^ w10725;
	assign w10707 = w10771 ^ w10705;
	assign w10766 = w10682 ^ w10707;
	assign w10713 = w10709 ^ w10707;
	assign w10681 = w10713 ^ w43819;
	assign w10718 = w46469 ^ w10713;
	assign w10768 = w10727 ^ w10718;
	assign w10764 = w10768 & w10767;
	assign w10763 = w10764 ^ w10766;
	assign w10762 = w10765 & w10763;
	assign w10670 = w10762 ^ w10718;
	assign w10724 = w46471 ^ w10681;
	assign w10759 = w10764 ^ w10724;
	assign w10758 = w10759 & w10760;
	assign w10677 = w10758 ^ w10722;
	assign w10756 = w10764 ^ w10758;
	assign w10755 = w10766 & w10756;
	assign w10676 = w10758 ^ w10775;
	assign w43824 = w10755 ^ w10773;
	assign w10747 = w43824 ^ w10725;
	assign w10745 = w10747 & w10784;
	assign w10736 = w10747 & w10788;
	assign w10714 = w46475 ^ w43824;
	assign w10754 = w10714 ^ w10677;
	assign w10735 = w10754 & w10785;
	assign w10744 = w10754 & w10783;
	assign w10757 = w10758 ^ w10766;
	assign w10734 = w10757 & w10789;
	assign w10671 = w10676 ^ w10772;
	assign w10753 = w10755 ^ w10763;
	assign w10743 = w10757 & w46476;
	assign w43823 = w10743 ^ w10745;
	assign w10673 = w10762 ^ w10774;
	assign w10669 = w10673 ^ w10709;
	assign w10668 = w46471 ^ w10669;
	assign w10672 = w46469 ^ w10669;
	assign w10749 = w10671 ^ w10672;
	assign w10730 = w10749 & w10792;
	assign w10739 = w10749 & w10781;
	assign w10761 = w10762 ^ w10724;
	assign w10731 = w10761 & w10787;
	assign w10740 = w10761 & w10780;
	assign w10752 = w10761 & w10753;
	assign w10717 = w10752 ^ w10727;
	assign w10748 = w10717 ^ w10670;
	assign w10733 = w10748 & w10793;
	assign w10751 = w10717 ^ w10719;
	assign w10741 = w10751 & w10790;
	assign w10732 = w10751 & w10786;
	assign w10684 = w10740 ^ w10741;
	assign w10675 = w10752 ^ w10776;
	assign w10702 = w10740 ^ w10732;
	assign w10742 = w10748 & w10778;
	assign w43822 = w10741 ^ w10742;
	assign w10667 = w10714 ^ w10675;
	assign w10674 = w10704 ^ w10667;
	assign w10700 = w10742 ^ w10733;
	assign w10746 = w10667 ^ w10668;
	assign w10729 = w10746 & w10794;
	assign w43821 = w10729 ^ w10730;
	assign w10698 = w10702 ^ w43821;
	assign w10701 = w43823 ^ w10698;
	assign w10798 = w10700 ^ w10701;
	assign w45214 = ~w10798;
	assign w9608 = w45836 ^ w45214;
	assign w10738 = w10746 & w10779;
	assign w10699 = w10738 ^ w10741;
	assign w10723 = w10738 ^ w43822;
	assign w10689 = w10734 ^ w10723;
	assign w10686 = ~w10689;
	assign w10683 = w10739 ^ w10723;
	assign w10696 = ~w10699;
	assign w10695 = w10738 ^ w10739;
	assign w10750 = w10671 ^ w10674;
	assign w10737 = w10750 & w10782;
	assign w10715 = w10733 ^ w10737;
	assign w10693 = ~w10715;
	assign w10697 = w10693 ^ w10698;
	assign w10797 = w10696 ^ w10697;
	assign w9657 = w45835 ^ w10797;
	assign w10692 = w10693 ^ w10731;
	assign w50689 = ~w10797;
	assign w10688 = w10692 ^ w43823;
	assign w10691 = w10730 ^ w10688;
	assign w10728 = w10750 & w10791;
	assign w10694 = w10739 ^ w10728;
	assign w23516 = w46459 ^ w23520;
	assign w23503 = w23520 & w23516;
	assign w46481 = w50322 ^ w451;
	assign w25979 = w46483 ^ w46481;
	assign w25981 = w46482 ^ w25979;
	assign w25956 = w46481 ^ w46482;
	assign w26057 = w46478 ^ w25981;
	assign w26054 = w46479 ^ w25981;
	assign w26056 = w25986 ^ w25981;
	assign w10690 = ~w10694;
	assign w10795 = w10690 ^ w10691;
	assign w50693 = ~w10795;
	assign w9652 = w45841 ^ w10795;
	assign w10711 = w10735 ^ w43821;
	assign w10687 = w10711 ^ w10688;
	assign w50690 = w10686 ^ w10687;
	assign w10712 = w10736 ^ w10711;
	assign w10716 = w10744 ^ w10712;
	assign w10685 = w10743 ^ w10716;
	assign w50691 = w10684 ^ w10685;
	assign w9604 = ~w50691;
	assign w9614 = w50697 ^ w9604;
	assign w10721 = w10745 ^ w10716;
	assign w50692 = w43822 ^ w10721;
	assign w9655 = w50698 ^ w50692;
	assign w10796 = w10721 ^ w10695;
	assign w50694 = ~w10796;
	assign w9650 = w45834 ^ w10796;
	assign w9611 = ~w50690;
	assign w9610 = w50696 ^ w9611;
	assign w50695 = w10712 ^ w10683;
	assign w9831 = w50695 ^ w50699;
	assign w9612 = ~w9831;
	assign w14208 = w46463 ^ w14165;
	assign w14243 = w14248 ^ w14208;
	assign w14242 = w14243 & w14244;
	assign w14160 = w14242 ^ w14259;
	assign w14240 = w14248 ^ w14242;
	assign w14239 = w14250 & w14240;
	assign w43968 = w14239 ^ w14257;
	assign w14198 = w46467 ^ w43968;
	assign w14231 = w43968 ^ w14209;
	assign w14241 = w14242 ^ w14250;
	assign w14227 = w14241 & w46468;
	assign w14218 = w14241 & w14273;
	assign w14220 = w14231 & w14272;
	assign w14155 = w14160 ^ w14256;
	assign w14233 = w14155 ^ w14156;
	assign w14214 = w14233 & w14276;
	assign w14223 = w14233 & w14265;
	assign w14229 = w14231 & w14268;
	assign w43967 = w14227 ^ w14229;
	assign w14237 = w14239 ^ w14247;
	assign w14245 = w14246 ^ w14208;
	assign w14215 = w14245 & w14271;
	assign w14236 = w14245 & w14237;
	assign w14201 = w14236 ^ w14211;
	assign w14232 = w14201 ^ w14154;
	assign w14217 = w14232 & w14277;
	assign w14235 = w14201 ^ w14203;
	assign w14225 = w14235 & w14274;
	assign w14216 = w14235 & w14270;
	assign w14224 = w14245 & w14264;
	assign w14168 = w14224 ^ w14225;
	assign w14186 = w14224 ^ w14216;
	assign w14159 = w14236 ^ w14260;
	assign w14151 = w14198 ^ w14159;
	assign w14230 = w14151 ^ w14152;
	assign w14213 = w14230 & w14278;
	assign w43537 = w14213 ^ w14214;
	assign w14182 = w14186 ^ w43537;
	assign w14158 = w14188 ^ w14151;
	assign w14234 = w14155 ^ w14158;
	assign w14212 = w14234 & w14275;
	assign w14178 = w14223 ^ w14212;
	assign w14174 = ~w14178;
	assign w14221 = w14234 & w14266;
	assign w14199 = w14217 ^ w14221;
	assign w14177 = ~w14199;
	assign w14176 = w14177 ^ w14215;
	assign w14172 = w14176 ^ w43967;
	assign w14175 = w14214 ^ w14172;
	assign w14279 = w14174 ^ w14175;
	assign w45282 = ~w14279;
	assign w9841 = w45282 ^ w45825;
	assign w9737 = w9841 ^ w50683;
	assign w14181 = w14177 ^ w14182;
	assign w14185 = w43967 ^ w14182;
	assign w14226 = w14232 & w14262;
	assign w14184 = w14226 ^ w14217;
	assign w14282 = w14184 ^ w14185;
	assign w45285 = ~w14282;
	assign w9863 = w45285 ^ w45820;
	assign w43966 = w14225 ^ w14226;
	assign w14222 = w14230 & w14263;
	assign w14179 = w14222 ^ w14223;
	assign w14183 = w14222 ^ w14225;
	assign w14180 = ~w14183;
	assign w14281 = w14180 ^ w14181;
	assign w14207 = w14222 ^ w43966;
	assign w14167 = w14223 ^ w14207;
	assign w14173 = w14218 ^ w14207;
	assign w14170 = ~w14173;
	assign w45284 = ~w14281;
	assign w9859 = w45284 ^ w45819;
	assign w14161 = w14242 ^ w14206;
	assign w14238 = w14198 ^ w14161;
	assign w14228 = w14238 & w14267;
	assign w14219 = w14238 & w14269;
	assign w14195 = w14219 ^ w43537;
	assign w14196 = w14220 ^ w14195;
	assign w50680 = w14196 ^ w14167;
	assign w9825 = w50680 ^ w50684;
	assign w9704 = w9825 ^ w45284;
	assign w14200 = w14228 ^ w14196;
	assign w14205 = w14229 ^ w14200;
	assign w50679 = w43966 ^ w14205;
	assign w9846 = w50679 ^ w50683;
	assign w14280 = w14205 ^ w14179;
	assign w9695 = ~w50679;
	assign w9694 = w9825 ^ w9695;
	assign w14171 = w14195 ^ w14172;
	assign w45283 = ~w14280;
	assign w9690 = w50680 ^ w45283;
	assign w50677 = w14170 ^ w14171;
	assign w9856 = w50677 ^ w50681;
	assign w9739 = w9856 ^ w45819;
	assign w14169 = w14227 ^ w14200;
	assign w50678 = w14168 ^ w14169;
	assign w9851 = w50678 ^ w50682;
	assign w9701 = w9825 ^ w50678;
	assign w15006 = w46605 ^ w15001;
	assign w15056 = w15015 ^ w15006;
	assign w15052 = w15056 & w15055;
	assign w15051 = w15052 ^ w15054;
	assign w15047 = w15052 ^ w15012;
	assign w15046 = w15047 & w15048;
	assign w15045 = w15046 ^ w15054;
	assign w15031 = w15045 & w46612;
	assign w15044 = w15052 ^ w15046;
	assign w15043 = w15054 & w15044;
	assign w15041 = w15043 ^ w15051;
	assign w43999 = w15043 ^ w15061;
	assign w15002 = w46611 ^ w43999;
	assign w14965 = w15046 ^ w15010;
	assign w15035 = w43999 ^ w15013;
	assign w15024 = w15035 & w15076;
	assign w15033 = w15035 & w15072;
	assign w15042 = w15002 ^ w14965;
	assign w15023 = w15042 & w15073;
	assign w15032 = w15042 & w15071;
	assign w44002 = w15031 ^ w15033;
	assign w15022 = w15045 & w15077;
	assign w15050 = w15053 & w15051;
	assign w14958 = w15050 ^ w15006;
	assign w14961 = w15050 ^ w15062;
	assign w15049 = w15050 ^ w15012;
	assign w15040 = w15049 & w15041;
	assign w15005 = w15040 ^ w15015;
	assign w15036 = w15005 ^ w14958;
	assign w15039 = w15005 ^ w15007;
	assign w15020 = w15039 & w15074;
	assign w15029 = w15039 & w15078;
	assign w15028 = w15049 & w15068;
	assign w14972 = w15028 ^ w15029;
	assign w15021 = w15036 & w15081;
	assign w15030 = w15036 & w15066;
	assign w14990 = w15028 ^ w15020;
	assign w44001 = w15029 ^ w15030;
	assign w14963 = w15040 ^ w15064;
	assign w14955 = w15002 ^ w14963;
	assign w14962 = w14992 ^ w14955;
	assign w14964 = w15046 ^ w15063;
	assign w14959 = w14964 ^ w15060;
	assign w15038 = w14959 ^ w14962;
	assign w15016 = w15038 & w15079;
	assign w14988 = w15030 ^ w15021;
	assign w14957 = w14961 ^ w14997;
	assign w14960 = w46605 ^ w14957;
	assign w15037 = w14959 ^ w14960;
	assign w15018 = w15037 & w15080;
	assign w15027 = w15037 & w15069;
	assign w14956 = w46607 ^ w14957;
	assign w15034 = w14955 ^ w14956;
	assign w15017 = w15034 & w15082;
	assign w43998 = w15017 ^ w15018;
	assign w14986 = w14990 ^ w43998;
	assign w14989 = w44002 ^ w14986;
	assign w14999 = w15023 ^ w43998;
	assign w15000 = w15024 ^ w14999;
	assign w15086 = w14988 ^ w14989;
	assign w14982 = w15027 ^ w15016;
	assign w14978 = ~w14982;
	assign w45302 = ~w15086;
	assign w15026 = w15034 & w15067;
	assign w15011 = w15026 ^ w44001;
	assign w14971 = w15027 ^ w15011;
	assign w14983 = w15026 ^ w15027;
	assign w14987 = w15026 ^ w15029;
	assign w14984 = ~w14987;
	assign w50507 = w15000 ^ w14971;
	assign w43085 = w50507 ^ w50519;
	assign w42884 = w43123 ^ w43085;
	assign w42839 = w43085 ^ w45302;
	assign w14977 = w15022 ^ w15011;
	assign w14974 = ~w14977;
	assign w15004 = w15032 ^ w15000;
	assign w15009 = w15033 ^ w15004;
	assign w15084 = w15009 ^ w14983;
	assign w50506 = ~w15084;
	assign w50505 = w44001 ^ w15009;
	assign w42879 = ~w50505;
	assign w43068 = w50518 ^ w42879;
	assign w14973 = w15031 ^ w15004;
	assign w50504 = w14972 ^ w14973;
	assign w43099 = w50504 ^ w50517;
	assign w43070 = w43099 ^ w43090;
	assign w43033 = w45963 ^ w50504;
	assign w15025 = w15038 & w15070;
	assign w15003 = w15021 ^ w15025;
	assign w14981 = ~w15003;
	assign w14985 = w14981 ^ w14986;
	assign w15085 = w14984 ^ w14985;
	assign w45309 = ~w15085;
	assign w42882 = w43091 ^ w45309;
	assign w15019 = w15049 & w15075;
	assign w14980 = w14981 ^ w15019;
	assign w14976 = w14980 ^ w44002;
	assign w14975 = w14999 ^ w14976;
	assign w14979 = w15018 ^ w14976;
	assign w15083 = w14978 ^ w14979;
	assign w45308 = ~w15083;
	assign w43108 = w45308 ^ w45664;
	assign w43066 = w43108 ^ w43096;
	assign w43052 = w15084 ^ w45308;
	assign w43042 = w43108 ^ w50514;
	assign w50503 = w14974 ^ w14975;
	assign w42841 = w43085 ^ w50503;
	assign w43161 = w42841 ^ w42842;
	assign w45965 = ~w43079;
	assign w42998 = w45965 ^ w50460;
	assign w50347 = w42997 ^ w42998;
	assign w46456 = w50347 ^ w476;
	assign w23436 = w46456 ^ w46454;
	assign w23522 = w46456 ^ w46453;
	assign w42911 = w45965 ^ w45584;
	assign w50326 = w42911 ^ w42912;
	assign w42874 = w45965 ^ w50462;
	assign w43147 = w42874 ^ w42875;
	assign w50346 = w43147 ^ w43144;
	assign w23518 = w23522 ^ w23450;
	assign w46457 = w50346 ^ w475;
	assign w23433 = w46459 ^ w46457;
	assign w23514 = w23433 ^ w23522;
	assign w23507 = w23514 & w23518;
	assign w23410 = w46457 ^ w46458;
	assign w23439 = w23507 ^ w23436;
	assign w23513 = w46460 ^ w23514;
	assign w23435 = w46458 ^ w23433;
	assign w23510 = w23440 ^ w23435;
	assign w23511 = w46454 ^ w23435;
	assign w23501 = w23522 & w23511;
	assign w23502 = w23517 & w23510;
	assign w23437 = w23501 ^ w23435;
	assign w23443 = w23439 ^ w23437;
	assign w23448 = w46453 ^ w23443;
	assign w23395 = w23436 ^ w46455;
	assign w23519 = w46460 ^ w23395;
	assign w23524 = w46458 ^ w46456;
	assign w23509 = w23434 ^ w23524;
	assign w23500 = w23524 & w23509;
	assign w23409 = w23500 ^ w23501;
	assign w23456 = w23409 ^ w23410;
	assign w23505 = w46460 & w23519;
	assign w23396 = w23436 ^ w23434;
	assign w23512 = w23433 ^ w23396;
	assign w23508 = w46455 ^ w23435;
	assign w23504 = w23523 & w23508;
	assign w23438 = w23504 ^ w23434;
	assign w23455 = w23456 ^ w23438;
	assign w23497 = w23503 ^ w23455;
	assign w46477 = w50326 ^ w455;
	assign w26067 = w46477 ^ w46482;
	assign w25980 = w46479 ^ w46477;
	assign w25942 = w25982 ^ w25980;
	assign w26058 = w25979 ^ w25942;
	assign w26068 = w46480 ^ w46477;
	assign w26047 = w26068 & w26057;
	assign w26064 = w26068 ^ w25996;
	assign w26060 = w25979 ^ w26068;
	assign w26045 = w26067 & w26058;
	assign w26055 = w25980 ^ w26070;
	assign w26069 = w46477 ^ w46483;
	assign w44457 = w26045 ^ w26051;
	assign w26050 = w26069 & w26054;
	assign w25984 = w26050 ^ w25980;
	assign w26059 = w46484 ^ w26060;
	assign w25983 = w26047 ^ w25981;
	assign w26053 = w26060 & w26064;
	assign w25985 = w26053 ^ w25982;
	assign w25989 = w25985 ^ w25983;
	assign w25957 = w25989 ^ w44457;
	assign w26000 = w46479 ^ w25957;
	assign w25994 = w46477 ^ w25989;
	assign w25995 = w44457 ^ w25980;
	assign w26063 = w25980 ^ w25986;
	assign w26048 = w26063 & w26056;
	assign w44458 = w26045 ^ w26048;
	assign w25958 = w25984 ^ w44458;
	assign w26042 = w25958 ^ w25983;
	assign w26061 = w25996 ^ w26063;
	assign w23499 = w23521 & w23512;
	assign w44351 = w23499 ^ w23505;
	assign w44352 = w23499 ^ w23502;
	assign w23412 = w23438 ^ w44352;
	assign w23496 = w23412 ^ w23437;
	assign w23449 = w44351 ^ w23434;
	assign w23452 = w23500 ^ w44352;
	assign w23408 = w23503 ^ w23452;
	assign w23490 = w46459 ^ w23408;
	assign w23411 = w23443 ^ w44351;
	assign w23454 = w46455 ^ w23411;
	assign w26052 = w26061 & w26059;
	assign w26046 = w26070 & w26055;
	assign w25998 = w26046 ^ w44458;
	assign w25954 = w26049 ^ w25998;
	assign w26036 = w46483 ^ w25954;
	assign w25955 = w26046 ^ w26047;
	assign w26002 = w25955 ^ w25956;
	assign w26003 = w26046 ^ w26052;
	assign w26041 = w26003 ^ w25995;
	assign w26044 = w26003 ^ w25994;
	assign w26001 = w26002 ^ w25984;
	assign w26043 = w26049 ^ w26001;
	assign w26040 = w26044 & w26043;
	assign w26039 = w26040 ^ w26042;
	assign w26035 = w26040 ^ w26000;
	assign w26034 = w26035 & w26036;
	assign w25953 = w26034 ^ w25998;
	assign w26032 = w26040 ^ w26034;
	assign w26031 = w26042 & w26032;
	assign w26029 = w26031 ^ w26039;
	assign w26033 = w26034 ^ w26042;
	assign w25952 = w26034 ^ w26051;
	assign w25947 = w25952 ^ w26048;
	assign w26010 = w26033 & w26065;
	assign w44461 = w26031 ^ w26049;
	assign w25990 = w46483 ^ w44461;
	assign w26030 = w25990 ^ w25953;
	assign w26011 = w26030 & w26061;
	assign w26020 = w26030 & w26059;
	assign w26023 = w44461 ^ w26001;
	assign w26021 = w26023 & w26060;
	assign w26012 = w26023 & w26064;
	assign w26019 = w26033 & w46484;
	assign w44460 = w26019 ^ w26021;
	assign w26038 = w26041 & w26039;
	assign w26037 = w26038 ^ w26000;
	assign w26028 = w26037 & w26029;
	assign w25951 = w26028 ^ w26052;
	assign w25993 = w26028 ^ w26003;
	assign w26027 = w25993 ^ w25995;
	assign w26017 = w26027 & w26066;
	assign w26016 = w26037 & w26056;
	assign w25960 = w26016 ^ w26017;
	assign w25949 = w26038 ^ w26050;
	assign w25945 = w25949 ^ w25985;
	assign w25948 = w46477 ^ w25945;
	assign w25943 = w25990 ^ w25951;
	assign w25950 = w25980 ^ w25943;
	assign w25944 = w46479 ^ w25945;
	assign w26022 = w25943 ^ w25944;
	assign w26014 = w26022 & w26055;
	assign w25975 = w26014 ^ w26017;
	assign w25972 = ~w25975;
	assign w26005 = w26022 & w26070;
	assign w26007 = w26037 & w26063;
	assign w26026 = w25947 ^ w25950;
	assign w26013 = w26026 & w26058;
	assign w26004 = w26026 & w26067;
	assign w26025 = w25947 ^ w25948;
	assign w26015 = w26025 & w26057;
	assign w25971 = w26014 ^ w26015;
	assign w25970 = w26015 ^ w26004;
	assign w25966 = ~w25970;
	assign w26008 = w26027 & w26062;
	assign w25978 = w26016 ^ w26008;
	assign w26006 = w26025 & w26068;
	assign w43572 = w26005 ^ w26006;
	assign w25974 = w25978 ^ w43572;
	assign w25977 = w44460 ^ w25974;
	assign w25987 = w26011 ^ w43572;
	assign w25988 = w26012 ^ w25987;
	assign w25992 = w26020 ^ w25988;
	assign w25961 = w26019 ^ w25992;
	assign w25997 = w26021 ^ w25992;
	assign w26072 = w25997 ^ w25971;
	assign w9814 = w50712 ^ w26072;
	assign w50707 = ~w26072;
	assign w9887 = w50707 ^ w45216;
	assign w50705 = w25960 ^ w25961;
	assign w25946 = w26038 ^ w25994;
	assign w26024 = w25993 ^ w25946;
	assign w26009 = w26024 & w26069;
	assign w25991 = w26009 ^ w26013;
	assign w25969 = ~w25991;
	assign w25973 = w25969 ^ w25974;
	assign w26073 = w25972 ^ w25973;
	assign w26018 = w26024 & w26054;
	assign w25976 = w26018 ^ w26009;
	assign w26074 = w25976 ^ w25977;
	assign w45576 = ~w26073;
	assign w9877 = w45576 ^ w45217;
	assign w9786 = ~w9877;
	assign w45577 = ~w26074;
	assign w9885 = w45577 ^ w45213;
	assign w44459 = w26017 ^ w26018;
	assign w25999 = w26014 ^ w44459;
	assign w25965 = w26010 ^ w25999;
	assign w25962 = ~w25965;
	assign w50706 = w44459 ^ w25997;
	assign w9628 = ~w50706;
	assign w9627 = w50710 ^ w9628;
	assign w9888 = w50706 ^ w50711;
	assign w25959 = w26015 ^ w25999;
	assign w50708 = w25988 ^ w25959;
	assign w9823 = w50708 ^ w50712;
	assign w23506 = w23515 & w23513;
	assign w23457 = w23500 ^ w23506;
	assign w23495 = w23457 ^ w23449;
	assign w23498 = w23457 ^ w23448;
	assign w23494 = w23498 & w23497;
	assign w23493 = w23494 ^ w23496;
	assign w23489 = w23494 ^ w23454;
	assign w23492 = w23495 & w23493;
	assign w23403 = w23492 ^ w23504;
	assign w23400 = w23492 ^ w23448;
	assign w23488 = w23489 & w23490;
	assign w23487 = w23488 ^ w23496;
	assign w23464 = w23487 & w23519;
	assign w23473 = w23487 & w46460;
	assign w23406 = w23488 ^ w23505;
	assign w23401 = w23406 ^ w23502;
	assign w23399 = w23403 ^ w23439;
	assign w23402 = w46453 ^ w23399;
	assign w23479 = w23401 ^ w23402;
	assign w23398 = w46455 ^ w23399;
	assign w23486 = w23494 ^ w23488;
	assign w23485 = w23496 & w23486;
	assign w23483 = w23485 ^ w23493;
	assign w23460 = w23479 & w23522;
	assign w23407 = w23488 ^ w23452;
	assign w23469 = w23479 & w23511;
	assign w44356 = w23485 ^ w23503;
	assign w23444 = w46459 ^ w44356;
	assign w23484 = w23444 ^ w23407;
	assign w23474 = w23484 & w23513;
	assign w23477 = w44356 ^ w23455;
	assign w23475 = w23477 & w23514;
	assign w44355 = w23473 ^ w23475;
	assign w23466 = w23477 & w23518;
	assign w23491 = w23492 ^ w23454;
	assign w23470 = w23491 & w23510;
	assign w23482 = w23491 & w23483;
	assign w23447 = w23482 ^ w23457;
	assign w23481 = w23447 ^ w23449;
	assign w23462 = w23481 & w23516;
	assign w23478 = w23447 ^ w23400;
	assign w23472 = w23478 & w23508;
	assign w23463 = w23478 & w23523;
	assign w23430 = w23472 ^ w23463;
	assign w23432 = w23470 ^ w23462;
	assign w23461 = w23491 & w23517;
	assign w23471 = w23481 & w23520;
	assign w23414 = w23470 ^ w23471;
	assign w44354 = w23471 ^ w23472;
	assign w23405 = w23482 ^ w23506;
	assign w23397 = w23444 ^ w23405;
	assign w23476 = w23397 ^ w23398;
	assign w23468 = w23476 & w23509;
	assign w23425 = w23468 ^ w23469;
	assign w23429 = w23468 ^ w23471;
	assign w23426 = ~w23429;
	assign w23453 = w23468 ^ w44354;
	assign w23419 = w23464 ^ w23453;
	assign w23416 = ~w23419;
	assign w23413 = w23469 ^ w23453;
	assign w23459 = w23476 & w23524;
	assign w44353 = w23459 ^ w23460;
	assign w23428 = w23432 ^ w44353;
	assign w23431 = w44355 ^ w23428;
	assign w23528 = w23430 ^ w23431;
	assign w23404 = w23434 ^ w23397;
	assign w23480 = w23401 ^ w23404;
	assign w23467 = w23480 & w23512;
	assign w23445 = w23463 ^ w23467;
	assign w23423 = ~w23445;
	assign w23427 = w23423 ^ w23428;
	assign w23527 = w23426 ^ w23427;
	assign w23422 = w23423 ^ w23461;
	assign w23418 = w23422 ^ w44355;
	assign w23458 = w23480 & w23521;
	assign w23424 = w23469 ^ w23458;
	assign w23420 = ~w23424;
	assign w45502 = ~w23527;
	assign w9891 = w45280 ^ w45502;
	assign w45503 = ~w23528;
	assign w9892 = w45281 ^ w45503;
	assign w23421 = w23460 ^ w23418;
	assign w23525 = w23420 ^ w23421;
	assign w45509 = ~w23525;
	assign w23465 = w23484 & w23515;
	assign w23441 = w23465 ^ w44353;
	assign w23417 = w23441 ^ w23418;
	assign w23442 = w23466 ^ w23441;
	assign w23446 = w23474 ^ w23442;
	assign w23415 = w23473 ^ w23446;
	assign w50664 = w23414 ^ w23415;
	assign w50667 = w23442 ^ w23413;
	assign w9836 = w50651 ^ w50667;
	assign w9578 = w9836 ^ w50649;
	assign w9732 = ~w9836;
	assign w50663 = w23416 ^ w23417;
	assign w9871 = w50648 ^ w50663;
	assign w9733 = ~w9871;
	assign w9761 = w9732 ^ w45502;
	assign w23451 = w23475 ^ w23446;
	assign w23526 = w23451 ^ w23425;
	assign w50666 = ~w23526;
	assign w50665 = w44354 ^ w23451;
	assign w45951 = ~w9823;
	assign w9811 = w45951 ^ w45576;
	assign w9626 = w45951 ^ w50705;
	assign w9895 = w9626 ^ w9627;
	assign w25968 = w25969 ^ w26007;
	assign w25964 = w25968 ^ w44460;
	assign w25963 = w25987 ^ w25964;
	assign w50704 = w25962 ^ w25963;
	assign w9862 = w50704 ^ w50709;
	assign w25967 = w26006 ^ w25964;
	assign w26071 = w25966 ^ w25967;
	assign w45575 = ~w26071;
	assign w9801 = w26072 ^ w45575;
	assign w45971 = ~w43421;
	assign w43323 = w45971 ^ w45586;
	assign w43321 = w43322 ^ w43323;
	assign w50159 = ~w43321;
	assign w46571 = w50159 ^ w1286;
	assign w10988 = w46571 ^ w46570;
	assign w11054 = w46571 ^ w11058;
	assign w43319 = w45971 ^ w50267;
	assign w50161 = w43318 ^ w43319;
	assign w46569 = w50161 ^ w1288;
	assign w10948 = w46569 ^ w46570;
	assign w43316 = w45971 ^ w50268;
	assign w50162 = w43315 ^ w43316;
	assign w11053 = w10988 ^ w11055;
	assign w46568 = w50162 ^ w1289;
	assign w11062 = w46570 ^ w46568;
	assign w10974 = w46568 ^ w46566;
	assign w10934 = w10974 ^ w10972;
	assign w11047 = w10972 ^ w11062;
	assign w11041 = w11058 & w11054;
	assign w10933 = w10974 ^ w46567;
	assign w11057 = w46572 ^ w10933;
	assign w11043 = w46572 & w11057;
	assign w11038 = w11062 & w11047;
	assign w10971 = w46571 ^ w46569;
	assign w10973 = w46570 ^ w10971;
	assign w11046 = w46567 ^ w10973;
	assign w11048 = w10978 ^ w10973;
	assign w11050 = w10971 ^ w10934;
	assign w11037 = w11059 & w11050;
	assign w11049 = w46566 ^ w10973;
	assign w43834 = w11037 ^ w11043;
	assign w10987 = w43834 ^ w10972;
	assign w11040 = w11055 & w11048;
	assign w43831 = w11037 ^ w11040;
	assign w10990 = w11038 ^ w43831;
	assign w10946 = w11041 ^ w10990;
	assign w11028 = w46571 ^ w10946;
	assign w11061 = w46565 ^ w46571;
	assign w11042 = w11061 & w11046;
	assign w11060 = w46568 ^ w46565;
	assign w11056 = w11060 ^ w10988;
	assign w11039 = w11060 & w11049;
	assign w10975 = w11039 ^ w10973;
	assign w10947 = w11038 ^ w11039;
	assign w11052 = w10971 ^ w11060;
	assign w11051 = w46572 ^ w11052;
	assign w11044 = w11053 & w11051;
	assign w11045 = w11052 & w11056;
	assign w10977 = w11045 ^ w10974;
	assign w10981 = w10977 ^ w10975;
	assign w10949 = w10981 ^ w43834;
	assign w10986 = w46565 ^ w10981;
	assign w10995 = w11038 ^ w11044;
	assign w11036 = w10995 ^ w10986;
	assign w10992 = w46567 ^ w10949;
	assign w10994 = w10947 ^ w10948;
	assign w11033 = w10995 ^ w10987;
	assign w10976 = w11042 ^ w10972;
	assign w10993 = w10994 ^ w10976;
	assign w11035 = w11041 ^ w10993;
	assign w10950 = w10976 ^ w43831;
	assign w11034 = w10950 ^ w10975;
	assign w11032 = w11036 & w11035;
	assign w11031 = w11032 ^ w11034;
	assign w11027 = w11032 ^ w10992;
	assign w11026 = w11027 & w11028;
	assign w11025 = w11026 ^ w11034;
	assign w11011 = w11025 & w46572;
	assign w11030 = w11033 & w11031;
	assign w11029 = w11030 ^ w10992;
	assign w11008 = w11029 & w11048;
	assign w10941 = w11030 ^ w11042;
	assign w11002 = w11025 & w11057;
	assign w10937 = w10941 ^ w10977;
	assign w10936 = w46567 ^ w10937;
	assign w10999 = w11029 & w11055;
	assign w10938 = w11030 ^ w10986;
	assign w10945 = w11026 ^ w10990;
	assign w10940 = w46565 ^ w10937;
	assign w11024 = w11032 ^ w11026;
	assign w11023 = w11034 & w11024;
	assign w11021 = w11023 ^ w11031;
	assign w11020 = w11029 & w11021;
	assign w10943 = w11020 ^ w11044;
	assign w10985 = w11020 ^ w10995;
	assign w11016 = w10985 ^ w10938;
	assign w11001 = w11016 & w11061;
	assign w43833 = w11023 ^ w11041;
	assign w10982 = w46571 ^ w43833;
	assign w11022 = w10982 ^ w10945;
	assign w11012 = w11022 & w11051;
	assign w11003 = w11022 & w11053;
	assign w11015 = w43833 ^ w10993;
	assign w11013 = w11015 & w11052;
	assign w43836 = w11011 ^ w11013;
	assign w11004 = w11015 & w11056;
	assign w11010 = w11016 & w11046;
	assign w10935 = w10982 ^ w10943;
	assign w10942 = w10972 ^ w10935;
	assign w11014 = w10935 ^ w10936;
	assign w11006 = w11014 & w11047;
	assign w10997 = w11014 & w11062;
	assign w11019 = w10985 ^ w10987;
	assign w11009 = w11019 & w11058;
	assign w10952 = w11008 ^ w11009;
	assign w43835 = w11009 ^ w11010;
	assign w11000 = w11019 & w11054;
	assign w10991 = w11006 ^ w43835;
	assign w10957 = w11002 ^ w10991;
	assign w10970 = w11008 ^ w11000;
	assign w10967 = w11006 ^ w11009;
	assign w10968 = w11010 ^ w11001;
	assign w10954 = ~w10957;
	assign w10964 = ~w10967;
	assign w10944 = w11026 ^ w11043;
	assign w10939 = w10944 ^ w11040;
	assign w11018 = w10939 ^ w10942;
	assign w11005 = w11018 & w11050;
	assign w10983 = w11001 ^ w11005;
	assign w10996 = w11018 & w11059;
	assign w10961 = ~w10983;
	assign w10960 = w10961 ^ w10999;
	assign w10956 = w10960 ^ w43836;
	assign w11017 = w10939 ^ w10940;
	assign w11007 = w11017 & w11049;
	assign w10963 = w11006 ^ w11007;
	assign w10951 = w11007 ^ w10991;
	assign w10962 = w11007 ^ w10996;
	assign w10958 = ~w10962;
	assign w10998 = w11017 & w11060;
	assign w10959 = w10998 ^ w10956;
	assign w11063 = w10958 ^ w10959;
	assign w45224 = ~w11063;
	assign w43098 = w45224 ^ w45579;
	assign w43069 = ~w43098;
	assign w43067 = w43069 ^ w45664;
	assign w50420 = w43067 ^ w43068;
	assign w43051 = w43096 ^ w45224;
	assign w43050 = w43051 ^ w43052;
	assign w50429 = ~w43050;
	assign w43030 = w43098 ^ w43090;
	assign w50444 = w45308 ^ w43030;
	assign w46374 = w50429 ^ w1355;
	assign w46383 = w50420 ^ w1346;
	assign w43832 = w10997 ^ w10998;
	assign w10966 = w10970 ^ w43832;
	assign w10969 = w43836 ^ w10966;
	assign w11066 = w10968 ^ w10969;
	assign w45219 = ~w11066;
	assign w43136 = w45302 ^ w45219;
	assign w43061 = w43136 ^ w43103;
	assign w43038 = w43136 ^ w43073;
	assign w50439 = w45574 ^ w43038;
	assign w50415 = w45219 ^ w42884;
	assign w42826 = w45574 ^ w45219;
	assign w46364 = w50439 ^ w1365;
	assign w46388 = w50415 ^ w1341;
	assign w10965 = w10961 ^ w10966;
	assign w11065 = w10964 ^ w10965;
	assign w45218 = ~w11065;
	assign w43128 = w45309 ^ w45218;
	assign w43059 = w43128 ^ w43091;
	assign w50425 = w50503 ^ w43059;
	assign w46378 = w50425 ^ w1351;
	assign w43047 = w45581 ^ w45218;
	assign w43037 = ~w43128;
	assign w43035 = w43037 ^ w43123;
	assign w50440 = w43035 ^ w43036;
	assign w46363 = w50440 ^ w1366;
	assign w42840 = w45659 ^ w45218;
	assign w43162 = w42839 ^ w42840;
	assign w50416 = w43162 ^ w43103;
	assign w46387 = w50416 ^ w1342;
	assign w10979 = w11003 ^ w43832;
	assign w10980 = w11004 ^ w10979;
	assign w10955 = w10979 ^ w10956;
	assign w10984 = w11012 ^ w10980;
	assign w10989 = w11013 ^ w10984;
	assign w50510 = w43835 ^ w10989;
	assign w43139 = w50505 ^ w50510;
	assign w50443 = w43145 ^ w43139;
	assign w43071 = w43085 ^ w50510;
	assign w50419 = w43070 ^ w43071;
	assign w46384 = w50419 ^ w1345;
	assign w43055 = w43139 ^ w43108;
	assign w50428 = w45579 ^ w43055;
	assign w43043 = w45224 ^ w50510;
	assign w50436 = w43042 ^ w43043;
	assign w46367 = w50436 ^ w1362;
	assign w11064 = w10989 ^ w10963;
	assign w46375 = w50428 ^ w1354;
	assign w45225 = ~w11064;
	assign w43138 = w50506 ^ w45225;
	assign w50421 = w45225 ^ w43066;
	assign w43049 = w43138 ^ w43073;
	assign w50430 = w50507 ^ w43049;
	assign w46373 = w50430 ^ w1356;
	assign w40854 = w46375 ^ w46373;
	assign w40941 = w46373 ^ w46378;
	assign w43041 = w43138 ^ w43098;
	assign w50437 = w45665 ^ w43041;
	assign w43040 = w45580 ^ w45225;
	assign w43028 = w43138 ^ w45664;
	assign w50445 = w43028 ^ w43029;
	assign w46358 = w50445 ^ w1371;
	assign w39922 = w46364 ^ w46358;
	assign w46366 = w50437 ^ w1363;
	assign w46382 = w50421 ^ w1347;
	assign w40052 = w46384 ^ w46382;
	assign w40056 = w46388 ^ w46382;
	assign w40136 = w46383 ^ w40056;
	assign w40132 = w46387 ^ w40136;
	assign w40011 = w40052 ^ w46383;
	assign w40135 = w46388 ^ w40011;
	assign w40121 = w46388 & w40135;
	assign w40119 = w40136 & w40132;
	assign w10953 = w11011 ^ w10984;
	assign w46359 = w50444 ^ w1370;
	assign w40002 = w46359 ^ w39922;
	assign w39998 = w46363 ^ w40002;
	assign w39985 = w40002 & w39998;
	assign w50511 = w10980 ^ w10951;
	assign w43074 = w50507 ^ w50511;
	assign w43088 = w50511 ^ w50515;
	assign w43065 = w50511 ^ w15084;
	assign w50422 = w43064 ^ w43065;
	assign w43063 = w43123 ^ w43074;
	assign w50423 = w45302 ^ w43063;
	assign w43048 = w43136 ^ w43088;
	assign w50431 = w45659 ^ w43048;
	assign w46372 = w50431 ^ w1357;
	assign w41664 = w46372 ^ w46366;
	assign w41744 = w46367 ^ w41664;
	assign w43045 = w43088 ^ w50518;
	assign w43039 = w43074 ^ w50519;
	assign w50438 = w43039 ^ w43040;
	assign w46365 = w50438 ^ w1364;
	assign w41658 = w46367 ^ w46365;
	assign w41741 = w41658 ^ w41664;
	assign w43027 = w43096 ^ w43074;
	assign w50446 = w50515 ^ w43027;
	assign w42827 = w43088 ^ w50512;
	assign w42825 = w43088 ^ w45658;
	assign w43168 = w42825 ^ w42826;
	assign w50432 = w43168 ^ w43128;
	assign w46357 = w50446 ^ w1372;
	assign w39916 = w46359 ^ w46357;
	assign w39999 = w39916 ^ w39922;
	assign w40005 = w46357 ^ w46363;
	assign w46371 = w50432 ^ w1358;
	assign w41740 = w46371 ^ w41744;
	assign w41747 = w46365 ^ w46371;
	assign w41727 = w41744 & w41740;
	assign w46380 = w50423 ^ w1349;
	assign w40860 = w46380 ^ w46374;
	assign w40937 = w40854 ^ w40860;
	assign w40940 = w46375 ^ w40860;
	assign w46381 = w50422 ^ w1348;
	assign w40050 = w46383 ^ w46381;
	assign w40138 = w46384 ^ w46381;
	assign w40133 = w40050 ^ w40056;
	assign w40012 = w40052 ^ w40050;
	assign w40139 = w46381 ^ w46387;
	assign w50509 = w10952 ^ w10953;
	assign w43093 = w50509 ^ w50513;
	assign w50418 = w43161 ^ w43093;
	assign w43044 = w43139 ^ w43093;
	assign w50435 = w43044 ^ w43045;
	assign w46368 = w50435 ^ w1361;
	assign w41660 = w46368 ^ w46366;
	assign w41746 = w46368 ^ w46365;
	assign w41620 = w41660 ^ w41658;
	assign w41619 = w41660 ^ w46367;
	assign w41743 = w46372 ^ w41619;
	assign w41729 = w46372 & w41743;
	assign w43032 = w43093 ^ w43091;
	assign w43031 = w43032 ^ w43033;
	assign w50442 = ~w43031;
	assign w46361 = w50442 ^ w1368;
	assign w39915 = w46363 ^ w46361;
	assign w42878 = w50509 ^ w42879;
	assign w46385 = w50418 ^ w1344;
	assign w40049 = w46387 ^ w46385;
	assign w40130 = w40049 ^ w40138;
	assign w40129 = w46388 ^ w40130;
	assign w40128 = w40049 ^ w40012;
	assign w46360 = w50443 ^ w1369;
	assign w39918 = w46360 ^ w46358;
	assign w40004 = w46360 ^ w46357;
	assign w39996 = w39915 ^ w40004;
	assign w39995 = w46364 ^ w39996;
	assign w39878 = w39918 ^ w39916;
	assign w39994 = w39915 ^ w39878;
	assign w39877 = w39918 ^ w46359;
	assign w40001 = w46364 ^ w39877;
	assign w39987 = w46364 & w40001;
	assign w50508 = w10954 ^ w10955;
	assign w43113 = w50503 ^ w50508;
	assign w43058 = w43113 ^ w43099;
	assign w43056 = ~w43058;
	assign w43046 = w43113 ^ w50516;
	assign w50433 = w43046 ^ w43047;
	assign w43034 = w43113 ^ w43103;
	assign w50441 = w50512 ^ w43034;
	assign w42883 = w45658 ^ w50508;
	assign w50417 = w42882 ^ w42883;
	assign w46386 = w50417 ^ w1343;
	assign w40051 = w46386 ^ w40049;
	assign w40127 = w46382 ^ w40051;
	assign w40124 = w46383 ^ w40051;
	assign w40126 = w40056 ^ w40051;
	assign w40066 = w46387 ^ w46386;
	assign w40131 = w40066 ^ w40133;
	assign w40134 = w40138 ^ w40066;
	assign w40140 = w46386 ^ w46384;
	assign w40125 = w40050 ^ w40140;
	assign w40026 = w46385 ^ w46386;
	assign w40137 = w46381 ^ w46386;
	assign w40123 = w40130 & w40134;
	assign w40055 = w40123 ^ w40052;
	assign w40122 = w40131 & w40129;
	assign w40120 = w40139 & w40124;
	assign w40054 = w40120 ^ w40050;
	assign w40118 = w40133 & w40126;
	assign w40117 = w40138 & w40127;
	assign w40053 = w40117 ^ w40051;
	assign w40059 = w40055 ^ w40053;
	assign w40064 = w46381 ^ w40059;
	assign w40116 = w40140 & w40125;
	assign w40073 = w40116 ^ w40122;
	assign w40114 = w40073 ^ w40064;
	assign w40025 = w40116 ^ w40117;
	assign w40072 = w40025 ^ w40026;
	assign w40071 = w40072 ^ w40054;
	assign w40113 = w40119 ^ w40071;
	assign w40115 = w40137 & w40128;
	assign w40110 = w40114 & w40113;
	assign w42828 = w50509 ^ w50508;
	assign w43167 = w42827 ^ w42828;
	assign w50434 = w43167 ^ w43099;
	assign w46369 = w50434 ^ w1360;
	assign w41657 = w46371 ^ w46369;
	assign w41738 = w41657 ^ w41746;
	assign w41737 = w46372 ^ w41738;
	assign w41736 = w41657 ^ w41620;
	assign w46362 = w50441 ^ w1367;
	assign w39917 = w46362 ^ w39915;
	assign w39993 = w46358 ^ w39917;
	assign w39990 = w46359 ^ w39917;
	assign w39992 = w39922 ^ w39917;
	assign w39932 = w46363 ^ w46362;
	assign w39997 = w39932 ^ w39999;
	assign w40000 = w40004 ^ w39932;
	assign w40006 = w46362 ^ w46360;
	assign w39991 = w39916 ^ w40006;
	assign w39892 = w46361 ^ w46362;
	assign w40003 = w46357 ^ w46362;
	assign w39989 = w39996 & w40000;
	assign w39921 = w39989 ^ w39918;
	assign w39988 = w39997 & w39995;
	assign w39986 = w40005 & w39990;
	assign w39920 = w39986 ^ w39916;
	assign w39984 = w39999 & w39992;
	assign w39983 = w40004 & w39993;
	assign w39919 = w39983 ^ w39917;
	assign w39925 = w39921 ^ w39919;
	assign w39930 = w46357 ^ w39925;
	assign w39982 = w40006 & w39991;
	assign w39939 = w39982 ^ w39988;
	assign w39980 = w39939 ^ w39930;
	assign w39891 = w39982 ^ w39983;
	assign w39938 = w39891 ^ w39892;
	assign w39937 = w39938 ^ w39920;
	assign w39979 = w39985 ^ w39937;
	assign w39981 = w40003 & w39994;
	assign w39976 = w39980 & w39979;
	assign w46370 = w50433 ^ w1359;
	assign w41659 = w46370 ^ w41657;
	assign w41735 = w46366 ^ w41659;
	assign w41732 = w46367 ^ w41659;
	assign w41734 = w41664 ^ w41659;
	assign w41674 = w46371 ^ w46370;
	assign w41739 = w41674 ^ w41741;
	assign w41742 = w41746 ^ w41674;
	assign w41748 = w46370 ^ w46368;
	assign w41733 = w41658 ^ w41748;
	assign w41634 = w46369 ^ w46370;
	assign w41745 = w46365 ^ w46370;
	assign w41731 = w41738 & w41742;
	assign w41663 = w41731 ^ w41660;
	assign w41730 = w41739 & w41737;
	assign w41728 = w41747 & w41732;
	assign w41662 = w41728 ^ w41658;
	assign w41726 = w41741 & w41734;
	assign w41725 = w41746 & w41735;
	assign w41661 = w41725 ^ w41659;
	assign w41667 = w41663 ^ w41661;
	assign w41672 = w46365 ^ w41667;
	assign w41724 = w41748 & w41733;
	assign w41681 = w41724 ^ w41730;
	assign w41722 = w41681 ^ w41672;
	assign w41633 = w41724 ^ w41725;
	assign w41680 = w41633 ^ w41634;
	assign w41679 = w41680 ^ w41662;
	assign w41721 = w41727 ^ w41679;
	assign w41723 = w41745 & w41736;
	assign w41718 = w41722 & w41721;
	assign w45044 = w39981 ^ w39987;
	assign w39931 = w45044 ^ w39916;
	assign w39977 = w39939 ^ w39931;
	assign w39893 = w39925 ^ w45044;
	assign w39936 = w46359 ^ w39893;
	assign w39971 = w39976 ^ w39936;
	assign w45045 = w39981 ^ w39984;
	assign w39934 = w39982 ^ w45045;
	assign w39890 = w39985 ^ w39934;
	assign w39972 = w46363 ^ w39890;
	assign w39970 = w39971 & w39972;
	assign w39968 = w39976 ^ w39970;
	assign w39889 = w39970 ^ w39934;
	assign w39888 = w39970 ^ w39987;
	assign w39883 = w39888 ^ w39984;
	assign w39894 = w39920 ^ w45045;
	assign w39978 = w39894 ^ w39919;
	assign w39969 = w39970 ^ w39978;
	assign w39975 = w39976 ^ w39978;
	assign w39974 = w39977 & w39975;
	assign w39973 = w39974 ^ w39936;
	assign w39885 = w39974 ^ w39986;
	assign w39881 = w39885 ^ w39921;
	assign w39884 = w46357 ^ w39881;
	assign w39961 = w39883 ^ w39884;
	assign w39882 = w39974 ^ w39930;
	assign w39880 = w46359 ^ w39881;
	assign w39967 = w39978 & w39968;
	assign w39965 = w39967 ^ w39975;
	assign w39964 = w39973 & w39965;
	assign w39929 = w39964 ^ w39939;
	assign w39963 = w39929 ^ w39931;
	assign w39887 = w39964 ^ w39988;
	assign w39960 = w39929 ^ w39882;
	assign w39955 = w39969 & w46364;
	assign w39954 = w39960 & w39990;
	assign w39953 = w39963 & w40002;
	assign w39952 = w39973 & w39992;
	assign w39896 = w39952 ^ w39953;
	assign w39951 = w39961 & w39993;
	assign w39946 = w39969 & w40001;
	assign w39945 = w39960 & w40005;
	assign w39912 = w39954 ^ w39945;
	assign w39944 = w39963 & w39998;
	assign w39914 = w39952 ^ w39944;
	assign w39943 = w39973 & w39999;
	assign w39942 = w39961 & w40004;
	assign w45046 = w39953 ^ w39954;
	assign w45048 = w39967 ^ w39985;
	assign w39926 = w46363 ^ w45048;
	assign w39966 = w39926 ^ w39889;
	assign w39879 = w39926 ^ w39887;
	assign w39886 = w39916 ^ w39879;
	assign w39962 = w39883 ^ w39886;
	assign w39958 = w39879 ^ w39880;
	assign w39956 = w39966 & w39995;
	assign w39950 = w39958 & w39991;
	assign w39911 = w39950 ^ w39953;
	assign w39908 = ~w39911;
	assign w39907 = w39950 ^ w39951;
	assign w39949 = w39962 & w39994;
	assign w39947 = w39966 & w39997;
	assign w39927 = w39945 ^ w39949;
	assign w39905 = ~w39927;
	assign w39904 = w39905 ^ w39943;
	assign w39941 = w39958 & w40006;
	assign w39940 = w39962 & w40003;
	assign w39906 = w39951 ^ w39940;
	assign w39902 = ~w39906;
	assign w43609 = w39941 ^ w39942;
	assign w39923 = w39947 ^ w43609;
	assign w39910 = w39914 ^ w43609;
	assign w39909 = w39905 ^ w39910;
	assign w40009 = w39908 ^ w39909;
	assign w39935 = w39950 ^ w45046;
	assign w39901 = w39946 ^ w39935;
	assign w39898 = ~w39901;
	assign w39895 = w39951 ^ w39935;
	assign w39959 = w45048 ^ w39937;
	assign w39957 = w39959 & w39996;
	assign w39948 = w39959 & w40000;
	assign w39924 = w39948 ^ w39923;
	assign w39928 = w39956 ^ w39924;
	assign w39933 = w39957 ^ w39928;
	assign w50719 = w45046 ^ w39933;
	assign w40008 = w39933 ^ w39907;
	assign w39897 = w39955 ^ w39928;
	assign w50718 = w39896 ^ w39897;
	assign w50720 = w39924 ^ w39895;
	assign w9848 = w50705 ^ w50718;
	assign w9807 = w9862 ^ w9848;
	assign w9805 = ~w9807;
	assign w45047 = w39955 ^ w39957;
	assign w39913 = w45047 ^ w39910;
	assign w40010 = w39912 ^ w39913;
	assign w39900 = w39904 ^ w45047;
	assign w39903 = w39942 ^ w39900;
	assign w40007 = w39902 ^ w39903;
	assign w39899 = w39923 ^ w39900;
	assign w50717 = w39898 ^ w39899;
	assign w9591 = w50718 ^ w50717;
	assign w9795 = w9862 ^ w50717;
	assign w45049 = w40115 ^ w40121;
	assign w40027 = w40059 ^ w45049;
	assign w40070 = w46383 ^ w40027;
	assign w40105 = w40110 ^ w40070;
	assign w40065 = w45049 ^ w40050;
	assign w40111 = w40073 ^ w40065;
	assign w45050 = w40115 ^ w40118;
	assign w40068 = w40116 ^ w45050;
	assign w40024 = w40119 ^ w40068;
	assign w40106 = w46387 ^ w40024;
	assign w40104 = w40105 & w40106;
	assign w40022 = w40104 ^ w40121;
	assign w40017 = w40022 ^ w40118;
	assign w40023 = w40104 ^ w40068;
	assign w40102 = w40110 ^ w40104;
	assign w40028 = w40054 ^ w45050;
	assign w40112 = w40028 ^ w40053;
	assign w40103 = w40104 ^ w40112;
	assign w40109 = w40110 ^ w40112;
	assign w40108 = w40111 & w40109;
	assign w40107 = w40108 ^ w40070;
	assign w40019 = w40108 ^ w40120;
	assign w40015 = w40019 ^ w40055;
	assign w40018 = w46381 ^ w40015;
	assign w40095 = w40017 ^ w40018;
	assign w40016 = w40108 ^ w40064;
	assign w40014 = w46383 ^ w40015;
	assign w40101 = w40112 & w40102;
	assign w40099 = w40101 ^ w40109;
	assign w40098 = w40107 & w40099;
	assign w40063 = w40098 ^ w40073;
	assign w40097 = w40063 ^ w40065;
	assign w40021 = w40098 ^ w40122;
	assign w40094 = w40063 ^ w40016;
	assign w40089 = w40103 & w46388;
	assign w40088 = w40094 & w40124;
	assign w40087 = w40097 & w40136;
	assign w40086 = w40107 & w40126;
	assign w40030 = w40086 ^ w40087;
	assign w40085 = w40095 & w40127;
	assign w40080 = w40103 & w40135;
	assign w40079 = w40094 & w40139;
	assign w40046 = w40088 ^ w40079;
	assign w40078 = w40097 & w40132;
	assign w40048 = w40086 ^ w40078;
	assign w40077 = w40107 & w40133;
	assign w40076 = w40095 & w40138;
	assign w45052 = w40087 ^ w40088;
	assign w45054 = w40101 ^ w40119;
	assign w40093 = w45054 ^ w40071;
	assign w40082 = w40093 & w40134;
	assign w40091 = w40093 & w40130;
	assign w45053 = w40089 ^ w40091;
	assign w40060 = w46387 ^ w45054;
	assign w40100 = w40060 ^ w40023;
	assign w40013 = w40060 ^ w40021;
	assign w40020 = w40050 ^ w40013;
	assign w40096 = w40017 ^ w40020;
	assign w40092 = w40013 ^ w40014;
	assign w40090 = w40100 & w40129;
	assign w40084 = w40092 & w40125;
	assign w40069 = w40084 ^ w45052;
	assign w40045 = w40084 ^ w40087;
	assign w40042 = ~w40045;
	assign w40041 = w40084 ^ w40085;
	assign w40035 = w40080 ^ w40069;
	assign w40032 = ~w40035;
	assign w40029 = w40085 ^ w40069;
	assign w40083 = w40096 & w40128;
	assign w40061 = w40079 ^ w40083;
	assign w40039 = ~w40061;
	assign w40038 = w40039 ^ w40077;
	assign w40034 = w40038 ^ w45053;
	assign w40037 = w40076 ^ w40034;
	assign w40081 = w40100 & w40131;
	assign w40075 = w40092 & w40140;
	assign w40074 = w40096 & w40137;
	assign w40040 = w40085 ^ w40074;
	assign w40036 = ~w40040;
	assign w40141 = w40036 ^ w40037;
	assign w45051 = w40075 ^ w40076;
	assign w40057 = w40081 ^ w45051;
	assign w40058 = w40082 ^ w40057;
	assign w40062 = w40090 ^ w40058;
	assign w40067 = w40091 ^ w40062;
	assign w50687 = w45052 ^ w40067;
	assign w40142 = w40067 ^ w40041;
	assign w40033 = w40057 ^ w40034;
	assign w50685 = w40032 ^ w40033;
	assign w40031 = w40089 ^ w40062;
	assign w50686 = w40030 ^ w40031;
	assign w9875 = w50686 ^ w50691;
	assign w50688 = w40058 ^ w40029;
	assign w9603 = w9604 ^ w50685;
	assign w9867 = w50687 ^ w50692;
	assign w9683 = w10795 ^ w50687;
	assign w9639 = ~w9867;
	assign w9827 = w50688 ^ w50695;
	assign w40044 = w40048 ^ w45051;
	assign w40047 = w45053 ^ w40044;
	assign w40144 = w40046 ^ w40047;
	assign w40043 = w40039 ^ w40044;
	assign w40143 = w40042 ^ w40043;
	assign w45116 = w41723 ^ w41729;
	assign w41635 = w41667 ^ w45116;
	assign w41678 = w46367 ^ w41635;
	assign w41713 = w41718 ^ w41678;
	assign w41673 = w45116 ^ w41658;
	assign w41719 = w41681 ^ w41673;
	assign w45117 = w41723 ^ w41726;
	assign w41676 = w41724 ^ w45117;
	assign w41632 = w41727 ^ w41676;
	assign w41714 = w46371 ^ w41632;
	assign w41712 = w41713 & w41714;
	assign w41631 = w41712 ^ w41676;
	assign w41630 = w41712 ^ w41729;
	assign w41625 = w41630 ^ w41726;
	assign w41710 = w41718 ^ w41712;
	assign w41636 = w41662 ^ w45117;
	assign w41720 = w41636 ^ w41661;
	assign w41711 = w41712 ^ w41720;
	assign w41717 = w41718 ^ w41720;
	assign w41716 = w41719 & w41717;
	assign w41715 = w41716 ^ w41678;
	assign w41627 = w41716 ^ w41728;
	assign w41623 = w41627 ^ w41663;
	assign w41626 = w46365 ^ w41623;
	assign w41703 = w41625 ^ w41626;
	assign w41624 = w41716 ^ w41672;
	assign w41622 = w46367 ^ w41623;
	assign w41709 = w41720 & w41710;
	assign w41707 = w41709 ^ w41717;
	assign w41706 = w41715 & w41707;
	assign w41671 = w41706 ^ w41681;
	assign w41705 = w41671 ^ w41673;
	assign w41629 = w41706 ^ w41730;
	assign w41702 = w41671 ^ w41624;
	assign w41697 = w41711 & w46372;
	assign w41696 = w41702 & w41732;
	assign w41695 = w41705 & w41744;
	assign w41694 = w41715 & w41734;
	assign w41638 = w41694 ^ w41695;
	assign w41693 = w41703 & w41735;
	assign w41688 = w41711 & w41743;
	assign w41687 = w41702 & w41747;
	assign w41654 = w41696 ^ w41687;
	assign w41686 = w41705 & w41740;
	assign w41656 = w41694 ^ w41686;
	assign w41685 = w41715 & w41741;
	assign w41684 = w41703 & w41746;
	assign w45119 = w41695 ^ w41696;
	assign w45121 = w41709 ^ w41727;
	assign w41701 = w45121 ^ w41679;
	assign w41699 = w41701 & w41738;
	assign w45120 = w41697 ^ w41699;
	assign w41690 = w41701 & w41742;
	assign w41668 = w46371 ^ w45121;
	assign w41708 = w41668 ^ w41631;
	assign w41621 = w41668 ^ w41629;
	assign w41628 = w41658 ^ w41621;
	assign w41704 = w41625 ^ w41628;
	assign w41700 = w41621 ^ w41622;
	assign w41698 = w41708 & w41737;
	assign w41692 = w41700 & w41733;
	assign w41677 = w41692 ^ w45119;
	assign w41653 = w41692 ^ w41695;
	assign w41650 = ~w41653;
	assign w41649 = w41692 ^ w41693;
	assign w41643 = w41688 ^ w41677;
	assign w41640 = ~w41643;
	assign w41637 = w41693 ^ w41677;
	assign w41691 = w41704 & w41736;
	assign w41669 = w41687 ^ w41691;
	assign w41647 = ~w41669;
	assign w41646 = w41647 ^ w41685;
	assign w41642 = w41646 ^ w45120;
	assign w41645 = w41684 ^ w41642;
	assign w41689 = w41708 & w41739;
	assign w41683 = w41700 & w41748;
	assign w41682 = w41704 & w41745;
	assign w41648 = w41693 ^ w41682;
	assign w41644 = ~w41648;
	assign w41749 = w41644 ^ w41645;
	assign w45118 = w41683 ^ w41684;
	assign w41665 = w41689 ^ w45118;
	assign w41641 = w41665 ^ w41642;
	assign w50659 = w41640 ^ w41641;
	assign w41666 = w41690 ^ w41665;
	assign w50662 = w41666 ^ w41637;
	assign w41670 = w41698 ^ w41666;
	assign w41639 = w41697 ^ w41670;
	assign w50660 = w41638 ^ w41639;
	assign w41675 = w41699 ^ w41670;
	assign w41750 = w41675 ^ w41649;
	assign w9828 = w50662 ^ w50667;
	assign w9625 = ~w50659;
	assign w9803 = w45280 ^ w9625;
	assign w9883 = w50660 ^ w50664;
	assign w9730 = w9883 ^ w9733;
	assign w50661 = w45119 ^ w41675;
	assign w9880 = w50661 ^ w50665;
	assign w41652 = w41656 ^ w45118;
	assign w41655 = w45120 ^ w41652;
	assign w41752 = w41654 ^ w41655;
	assign w41651 = w41647 ^ w41652;
	assign w41751 = w41650 ^ w41651;
	assign w50658 = ~w41751;
	assign w9750 = w45502 ^ w41751;
	assign w9618 = w41751 ^ w45281;
	assign w9834 = w50708 ^ w50720;
	assign w9588 = w9834 ^ w45577;
	assign w9590 = w9834 ^ w50704;
	assign w9910 = w9590 ^ w9591;
	assign w9621 = w9828 ^ w45503;
	assign w9606 = w50692 ^ w50686;
	assign w9642 = ~w9875;
	assign w9624 = w50660 ^ w9625;
	assign w9820 = w9834 ^ w50711;
	assign w9817 = w50719 ^ w9628;
	assign w45826 = ~w40008;
	assign w45827 = ~w40009;
	assign w9632 = w45827 ^ w50709;
	assign w45828 = ~w40010;
	assign w9589 = w45828 ^ w45217;
	assign w9911 = w9588 ^ w9589;
	assign w45830 = ~w40142;
	assign w9675 = w50695 ^ w45830;
	assign w9853 = w45830 ^ w50694;
	assign w45831 = ~w40143;
	assign w9889 = w45831 ^ w50689;
	assign w9686 = w9611 ^ w45831;
	assign w45832 = ~w40144;
	assign w9890 = w45832 ^ w45214;
	assign w9659 = w9890 ^ w9831;
	assign w9600 = w10797 ^ w45832;
	assign w45833 = ~w40007;
	assign w9777 = w9887 ^ w45833;
	assign w9857 = w45575 ^ w45833;
	assign w9804 = w9888 ^ w9857;
	assign w45837 = ~w40141;
	assign w9678 = w10796 ^ w45837;
	assign w9860 = w45837 ^ w50693;
	assign w45862 = ~w41749;
	assign w9876 = w45862 ^ w45509;
	assign w9699 = w9876 ^ w50650;
	assign w9697 = ~w9699;
	assign w45863 = ~w41750;
	assign w9873 = w45863 ^ w50666;
	assign w9680 = w9873 ^ w45278;
	assign w45864 = ~w41752;
	assign w9622 = w45280 ^ w45864;
	assign w9897 = w9621 ^ w9622;
	assign w45895 = ~w9827;
	assign w9672 = w45895 ^ w45831;
	assign w9666 = w45895 ^ w50687;
	assign w9668 = w45895 ^ w50686;
	assign w9788 = w9823 ^ w50720;
	assign w45954 = ~w9828;
	assign w9660 = w45954 ^ w45279;
	assign w9623 = w45954 ^ w50663;
	assign w9896 = w9623 ^ w9624;
	assign w9747 = w45954 ^ w50661;
	assign w45962 = ~w43074;
	assign w43062 = w45962 ^ w45309;
	assign w43060 = w43061 ^ w43062;
	assign w50424 = ~w43060;
	assign w46379 = w50424 ^ w1350;
	assign w40936 = w46379 ^ w40940;
	assign w40870 = w46379 ^ w46378;
	assign w40935 = w40870 ^ w40937;
	assign w40943 = w46373 ^ w46379;
	assign w40923 = w40940 & w40936;
	assign w43057 = w45962 ^ w50513;
	assign w50426 = w43056 ^ w43057;
	assign w42877 = w45962 ^ w50504;
	assign w43146 = w42877 ^ w42878;
	assign w50427 = w43146 ^ w43090;
	assign w46376 = w50427 ^ w1353;
	assign w40856 = w46376 ^ w46374;
	assign w40942 = w46376 ^ w46373;
	assign w40938 = w40942 ^ w40870;
	assign w40944 = w46378 ^ w46376;
	assign w40929 = w40854 ^ w40944;
	assign w40816 = w40856 ^ w40854;
	assign w40815 = w40856 ^ w46375;
	assign w40939 = w46380 ^ w40815;
	assign w40925 = w46380 & w40939;
	assign w40920 = w40944 & w40929;
	assign w46377 = w50426 ^ w1352;
	assign w40853 = w46379 ^ w46377;
	assign w40855 = w46378 ^ w40853;
	assign w40931 = w46374 ^ w40855;
	assign w40928 = w46375 ^ w40855;
	assign w40930 = w40860 ^ w40855;
	assign w40934 = w40853 ^ w40942;
	assign w40933 = w46380 ^ w40934;
	assign w40830 = w46377 ^ w46378;
	assign w40932 = w40853 ^ w40816;
	assign w40927 = w40934 & w40938;
	assign w40859 = w40927 ^ w40856;
	assign w40926 = w40935 & w40933;
	assign w40877 = w40920 ^ w40926;
	assign w40924 = w40943 & w40928;
	assign w40858 = w40924 ^ w40854;
	assign w40922 = w40937 & w40930;
	assign w40921 = w40942 & w40931;
	assign w40857 = w40921 ^ w40855;
	assign w40863 = w40859 ^ w40857;
	assign w40868 = w46373 ^ w40863;
	assign w40918 = w40877 ^ w40868;
	assign w40829 = w40920 ^ w40921;
	assign w40876 = w40829 ^ w40830;
	assign w40875 = w40876 ^ w40858;
	assign w40917 = w40923 ^ w40875;
	assign w40919 = w40941 & w40932;
	assign w40914 = w40918 & w40917;
	assign w45083 = w40919 ^ w40925;
	assign w40831 = w40863 ^ w45083;
	assign w40874 = w46375 ^ w40831;
	assign w40909 = w40914 ^ w40874;
	assign w40869 = w45083 ^ w40854;
	assign w40915 = w40877 ^ w40869;
	assign w45084 = w40919 ^ w40922;
	assign w40872 = w40920 ^ w45084;
	assign w40828 = w40923 ^ w40872;
	assign w40910 = w46379 ^ w40828;
	assign w40908 = w40909 & w40910;
	assign w40827 = w40908 ^ w40872;
	assign w40906 = w40914 ^ w40908;
	assign w40826 = w40908 ^ w40925;
	assign w40821 = w40826 ^ w40922;
	assign w40832 = w40858 ^ w45084;
	assign w40916 = w40832 ^ w40857;
	assign w40907 = w40908 ^ w40916;
	assign w40913 = w40914 ^ w40916;
	assign w40912 = w40915 & w40913;
	assign w40911 = w40912 ^ w40874;
	assign w40823 = w40912 ^ w40924;
	assign w40819 = w40823 ^ w40859;
	assign w40822 = w46373 ^ w40819;
	assign w40899 = w40821 ^ w40822;
	assign w40820 = w40912 ^ w40868;
	assign w40818 = w46375 ^ w40819;
	assign w40905 = w40916 & w40906;
	assign w40903 = w40905 ^ w40913;
	assign w40902 = w40911 & w40903;
	assign w40867 = w40902 ^ w40877;
	assign w40901 = w40867 ^ w40869;
	assign w40825 = w40902 ^ w40926;
	assign w40898 = w40867 ^ w40820;
	assign w40893 = w40907 & w46380;
	assign w40892 = w40898 & w40928;
	assign w40891 = w40901 & w40940;
	assign w40890 = w40911 & w40930;
	assign w40834 = w40890 ^ w40891;
	assign w40889 = w40899 & w40931;
	assign w40884 = w40907 & w40939;
	assign w40883 = w40898 & w40943;
	assign w40850 = w40892 ^ w40883;
	assign w40882 = w40901 & w40936;
	assign w40852 = w40890 ^ w40882;
	assign w40881 = w40911 & w40937;
	assign w40880 = w40899 & w40942;
	assign w45086 = w40891 ^ w40892;
	assign w45088 = w40905 ^ w40923;
	assign w40897 = w45088 ^ w40875;
	assign w40895 = w40897 & w40934;
	assign w45087 = w40893 ^ w40895;
	assign w40886 = w40897 & w40938;
	assign w40864 = w46379 ^ w45088;
	assign w40904 = w40864 ^ w40827;
	assign w40817 = w40864 ^ w40825;
	assign w40824 = w40854 ^ w40817;
	assign w40900 = w40821 ^ w40824;
	assign w40896 = w40817 ^ w40818;
	assign w40894 = w40904 & w40933;
	assign w40888 = w40896 & w40929;
	assign w40873 = w40888 ^ w45086;
	assign w40849 = w40888 ^ w40891;
	assign w40846 = ~w40849;
	assign w40845 = w40888 ^ w40889;
	assign w40839 = w40884 ^ w40873;
	assign w40836 = ~w40839;
	assign w40833 = w40889 ^ w40873;
	assign w40887 = w40900 & w40932;
	assign w40865 = w40883 ^ w40887;
	assign w40843 = ~w40865;
	assign w40842 = w40843 ^ w40881;
	assign w40838 = w40842 ^ w45087;
	assign w40841 = w40880 ^ w40838;
	assign w40885 = w40904 & w40935;
	assign w40879 = w40896 & w40944;
	assign w40878 = w40900 & w40941;
	assign w40844 = w40889 ^ w40878;
	assign w40840 = ~w40844;
	assign w40945 = w40840 ^ w40841;
	assign w45085 = w40879 ^ w40880;
	assign w40861 = w40885 ^ w45085;
	assign w40837 = w40861 ^ w40838;
	assign w50673 = w40836 ^ w40837;
	assign w40862 = w40886 ^ w40861;
	assign w50676 = w40862 ^ w40833;
	assign w40866 = w40894 ^ w40862;
	assign w40835 = w40893 ^ w40866;
	assign w50674 = w40834 ^ w40835;
	assign w40871 = w40895 ^ w40866;
	assign w40946 = w40871 ^ w40845;
	assign w9585 = ~w50674;
	assign w9597 = w50678 ^ w9585;
	assign w9833 = w50676 ^ w50680;
	assign w9598 = ~w9833;
	assign w9596 = w9598 ^ w50683;
	assign w9907 = w9596 ^ w9597;
	assign w9594 = w9833 ^ w50682;
	assign w9592 = w9833 ^ w45819;
	assign w50675 = w45086 ^ w40871;
	assign w40848 = w40852 ^ w45085;
	assign w40851 = w45087 ^ w40848;
	assign w40948 = w40850 ^ w40851;
	assign w40847 = w40843 ^ w40848;
	assign w40947 = w40846 ^ w40847;
	assign w50672 = ~w40947;
	assign w9713 = w45284 ^ w40947;
	assign w9710 = w9695 ^ w50675;
	assign w9595 = w50677 ^ w50673;
	assign w9908 = w9594 ^ w9595;
	assign w45842 = ~w40948;
	assign w9593 = w45285 ^ w45842;
	assign w9909 = w9592 ^ w9593;
	assign w45848 = ~w40945;
	assign w45849 = ~w40946;
	assign w9716 = w9825 ^ w45849;
	assign w9708 = w45849 ^ w45848;
	assign w9843 = w45849 ^ w45283;
	assign w9691 = w9843 ^ w9841;
	assign w9735 = w9843 ^ w45818;
	assign w9882 = w50685 ^ w50690;
	assign w9658 = ~w9882;
	assign w45972 = ~w43419;
	assign w43241 = w45972 ^ w45314;
	assign w50207 = w43240 ^ w43241;
	assign w46523 = w50207 ^ w1270;
	assign w29278 = w46523 ^ w29282;
	assign w43236 = w45972 ^ w50295;
	assign w50209 = w43235 ^ w43236;
	assign w43233 = w45972 ^ w50296;
	assign w50210 = w43232 ^ w43233;
	assign w46520 = w50210 ^ w1273;
	assign w29198 = w46520 ^ w46518;
	assign w29158 = w29198 ^ w29196;
	assign w29285 = w46517 ^ w46523;
	assign w29284 = w46520 ^ w46517;
	assign w29265 = w29282 & w29278;
	assign w29286 = w46522 ^ w46520;
	assign w29271 = w29196 ^ w29286;
	assign w46521 = w50209 ^ w1272;
	assign w29172 = w46521 ^ w46522;
	assign w29195 = w46523 ^ w46521;
	assign w29276 = w29195 ^ w29284;
	assign w29274 = w29195 ^ w29158;
	assign w29275 = w46524 ^ w29276;
	assign w29261 = w29283 & w29274;
	assign w29197 = w46522 ^ w29195;
	assign w29273 = w46518 ^ w29197;
	assign w29270 = w46519 ^ w29197;
	assign w29272 = w29202 ^ w29197;
	assign w29264 = w29279 & w29272;
	assign w29263 = w29284 & w29273;
	assign w29199 = w29263 ^ w29197;
	assign w29262 = w29286 & w29271;
	assign w44592 = w29261 ^ w29264;
	assign w29214 = w29262 ^ w44592;
	assign w29170 = w29265 ^ w29214;
	assign w29252 = w46523 ^ w29170;
	assign w29171 = w29262 ^ w29263;
	assign w29218 = w29171 ^ w29172;
	assign w29266 = w29285 & w29270;
	assign w29200 = w29266 ^ w29196;
	assign w29174 = w29200 ^ w44592;
	assign w29258 = w29174 ^ w29199;
	assign w29217 = w29218 ^ w29200;
	assign w29259 = w29265 ^ w29217;
	assign w29157 = w29198 ^ w46519;
	assign w29281 = w46524 ^ w29157;
	assign w29267 = w46524 & w29281;
	assign w44595 = w29261 ^ w29267;
	assign w29211 = w44595 ^ w29196;
	assign w29212 = w46523 ^ w46522;
	assign w29280 = w29284 ^ w29212;
	assign w29269 = w29276 & w29280;
	assign w29277 = w29212 ^ w29279;
	assign w29268 = w29277 & w29275;
	assign w29201 = w29269 ^ w29198;
	assign w29205 = w29201 ^ w29199;
	assign w29210 = w46517 ^ w29205;
	assign w29173 = w29205 ^ w44595;
	assign w29216 = w46519 ^ w29173;
	assign w29219 = w29262 ^ w29268;
	assign w29260 = w29219 ^ w29210;
	assign w29256 = w29260 & w29259;
	assign w29251 = w29256 ^ w29216;
	assign w29250 = w29251 & w29252;
	assign w29248 = w29256 ^ w29250;
	assign w29247 = w29258 & w29248;
	assign w29249 = w29250 ^ w29258;
	assign w29226 = w29249 & w29281;
	assign w29235 = w29249 & w46524;
	assign w29168 = w29250 ^ w29267;
	assign w44594 = w29247 ^ w29265;
	assign w29239 = w44594 ^ w29217;
	assign w29228 = w29239 & w29280;
	assign w29237 = w29239 & w29276;
	assign w29206 = w46523 ^ w44594;
	assign w29163 = w29168 ^ w29264;
	assign w44597 = w29235 ^ w29237;
	assign w29169 = w29250 ^ w29214;
	assign w29246 = w29206 ^ w29169;
	assign w29227 = w29246 & w29277;
	assign w29236 = w29246 & w29275;
	assign w29255 = w29256 ^ w29258;
	assign w29245 = w29247 ^ w29255;
	assign w29257 = w29219 ^ w29211;
	assign w29254 = w29257 & w29255;
	assign w29165 = w29254 ^ w29266;
	assign w29161 = w29165 ^ w29201;
	assign w29164 = w46517 ^ w29161;
	assign w29253 = w29254 ^ w29216;
	assign w29232 = w29253 & w29272;
	assign w29244 = w29253 & w29245;
	assign w29209 = w29244 ^ w29219;
	assign w29243 = w29209 ^ w29211;
	assign w29167 = w29244 ^ w29268;
	assign w29159 = w29206 ^ w29167;
	assign w29166 = w29196 ^ w29159;
	assign w29233 = w29243 & w29282;
	assign w29176 = w29232 ^ w29233;
	assign w29242 = w29163 ^ w29166;
	assign w29220 = w29242 & w29283;
	assign w29229 = w29242 & w29274;
	assign w29162 = w29254 ^ w29210;
	assign w29223 = w29253 & w29279;
	assign w29241 = w29163 ^ w29164;
	assign w29231 = w29241 & w29273;
	assign w29186 = w29231 ^ w29220;
	assign w29222 = w29241 & w29284;
	assign w29182 = ~w29186;
	assign w29160 = w46519 ^ w29161;
	assign w29238 = w29159 ^ w29160;
	assign w29221 = w29238 & w29286;
	assign w29230 = w29238 & w29271;
	assign w29187 = w29230 ^ w29231;
	assign w29191 = w29230 ^ w29233;
	assign w29188 = ~w29191;
	assign w44593 = w29221 ^ w29222;
	assign w29203 = w29227 ^ w44593;
	assign w29204 = w29228 ^ w29203;
	assign w29208 = w29236 ^ w29204;
	assign w29213 = w29237 ^ w29208;
	assign w29177 = w29235 ^ w29208;
	assign w50500 = w29176 ^ w29177;
	assign w43115 = w50496 ^ w50500;
	assign w42918 = w42909 ^ w43115;
	assign w50394 = w42918 ^ w42919;
	assign w42888 = w42890 ^ w43115;
	assign w42860 = w42863 ^ w50500;
	assign w43153 = w42860 ^ w42861;
	assign w50402 = w43153 ^ w43126;
	assign w46409 = w50394 ^ w395;
	assign w46401 = w50402 ^ w403;
	assign w29288 = w29213 ^ w29187;
	assign w29240 = w29209 ^ w29162;
	assign w29234 = w29240 & w29270;
	assign w44596 = w29233 ^ w29234;
	assign w50501 = w44596 ^ w29213;
	assign w42864 = w42863 ^ w50501;
	assign w43152 = w42864 ^ w42865;
	assign w50403 = w43152 ^ w43118;
	assign w46400 = w50403 ^ w404;
	assign w43106 = w50497 ^ w50501;
	assign w42887 = w43111 ^ w43106;
	assign w50412 = w45299 ^ w42887;
	assign w42916 = w42893 ^ w43106;
	assign w50395 = w42916 ^ w42917;
	assign w46408 = w50395 ^ w396;
	assign w29215 = w29230 ^ w44596;
	assign w29181 = w29226 ^ w29215;
	assign w29178 = ~w29181;
	assign w29225 = w29240 & w29285;
	assign w29207 = w29225 ^ w29229;
	assign w29192 = w29234 ^ w29225;
	assign w29185 = ~w29207;
	assign w29184 = w29185 ^ w29223;
	assign w29180 = w29184 ^ w44597;
	assign w29179 = w29203 ^ w29180;
	assign w50499 = w29178 ^ w29179;
	assign w43125 = w50495 ^ w50499;
	assign w42938 = ~w43125;
	assign w42920 = w43140 ^ w43125;
	assign w50393 = w50484 ^ w42920;
	assign w42907 = w42909 ^ w50499;
	assign w50401 = w42907 ^ w42908;
	assign w42891 = w42893 ^ w43125;
	assign w46410 = w50393 ^ w394;
	assign w42820 = w46410 ^ w46408;
	assign w42706 = w46409 ^ w46410;
	assign w29183 = w29222 ^ w29180;
	assign w29287 = w29182 ^ w29183;
	assign w46402 = w50401 ^ w402;
	assign w41882 = w46402 ^ w46400;
	assign w41768 = w46401 ^ w46402;
	assign w29175 = w29231 ^ w29215;
	assign w50502 = w29204 ^ w29175;
	assign w43075 = w50498 ^ w50502;
	assign w43083 = w50487 ^ w50502;
	assign w42913 = w43104 ^ w43075;
	assign w50398 = w50487 ^ w42913;
	assign w46405 = w50398 ^ w399;
	assign w42818 = w46408 ^ w46405;
	assign w42817 = w46405 ^ w46410;
	assign w42900 = w45899 ^ w50502;
	assign w50406 = w42900 ^ w42901;
	assign w42899 = w43141 ^ w43075;
	assign w50407 = w45294 ^ w42899;
	assign w46396 = w50407 ^ w408;
	assign w42856 = w43083 ^ w50500;
	assign w43155 = w42856 ^ w42857;
	assign w50387 = w43155 ^ w43106;
	assign w46416 = w50387 ^ w388;
	assign w42852 = ~w43083;
	assign w42853 = w42852 ^ w50499;
	assign w43156 = w42853 ^ w42854;
	assign w50386 = w43156 ^ w43115;
	assign w46397 = w50406 ^ w407;
	assign w41880 = w46400 ^ w46397;
	assign w41879 = w46397 ^ w46402;
	assign w46417 = w50386 ^ w387;
	assign w46391 = w50412 ^ w413;
	assign w45668 = ~w29287;
	assign w43100 = w45299 ^ w45668;
	assign w42935 = w43100 ^ w50501;
	assign w42933 = ~w42935;
	assign w50388 = w42933 ^ w42934;
	assign w42915 = w43118 ^ w43100;
	assign w50396 = w45291 ^ w42915;
	assign w42905 = w43111 ^ w45668;
	assign w50404 = w42905 ^ w42906;
	assign w42886 = w43104 ^ w43100;
	assign w50413 = w45300 ^ w42886;
	assign w46407 = w50396 ^ w397;
	assign w42730 = w46407 ^ w46405;
	assign w42805 = w42730 ^ w42820;
	assign w42796 = w42820 & w42805;
	assign w46415 = w50388 ^ w389;
	assign w46390 = w50413 ^ w414;
	assign w39386 = w46396 ^ w46390;
	assign w39466 = w46391 ^ w39386;
	assign w46399 = w50404 ^ w405;
	assign w41792 = w46399 ^ w46397;
	assign w41867 = w41792 ^ w41882;
	assign w41858 = w41882 & w41867;
	assign w45669 = ~w29288;
	assign w43089 = w45300 ^ w45669;
	assign w42928 = w43089 ^ w45668;
	assign w42927 = w42928 ^ w42929;
	assign w50389 = ~w42927;
	assign w42925 = w43075 ^ w45669;
	assign w50390 = w42925 ^ w42926;
	assign w42914 = w43111 ^ w43089;
	assign w50397 = w45292 ^ w42914;
	assign w46406 = w50397 ^ w398;
	assign w42732 = w46408 ^ w46406;
	assign w42692 = w42732 ^ w42730;
	assign w42691 = w42732 ^ w46407;
	assign w42904 = w43104 ^ w45669;
	assign w42902 = ~w42904;
	assign w50405 = w42902 ^ w42903;
	assign w42885 = w43089 ^ w43078;
	assign w50414 = w50498 ^ w42885;
	assign w46398 = w50405 ^ w406;
	assign w41794 = w46400 ^ w46398;
	assign w41754 = w41794 ^ w41792;
	assign w41753 = w41794 ^ w46399;
	assign w46389 = w50414 ^ w415;
	assign w39380 = w46391 ^ w46389;
	assign w39463 = w39380 ^ w39386;
	assign w46413 = w50390 ^ w391;
	assign w41926 = w46415 ^ w46413;
	assign w42014 = w46416 ^ w46413;
	assign w46414 = w50389 ^ w390;
	assign w41928 = w46416 ^ w46414;
	assign w41888 = w41928 ^ w41926;
	assign w41887 = w41928 ^ w46415;
	assign w29224 = w29243 & w29278;
	assign w29194 = w29232 ^ w29224;
	assign w29190 = w29194 ^ w44593;
	assign w29189 = w29185 ^ w29190;
	assign w29289 = w29188 ^ w29189;
	assign w29193 = w44597 ^ w29190;
	assign w29290 = w29192 ^ w29193;
	assign w45662 = ~w29289;
	assign w43129 = w45301 ^ w45662;
	assign w42936 = w42938 ^ w45662;
	assign w50385 = w42936 ^ w42937;
	assign w42922 = w43141 ^ w43129;
	assign w42921 = w42922 ^ w42923;
	assign w50392 = ~w42921;
	assign w46411 = w50392 ^ w393;
	assign w42729 = w46411 ^ w46409;
	assign w42731 = w46410 ^ w42729;
	assign w42807 = w46406 ^ w42731;
	assign w42804 = w46407 ^ w42731;
	assign w42810 = w42729 ^ w42818;
	assign w42746 = w46411 ^ w46410;
	assign w42814 = w42818 ^ w42746;
	assign w42808 = w42729 ^ w42692;
	assign w42819 = w46405 ^ w46411;
	assign w42803 = w42810 & w42814;
	assign w42735 = w42803 ^ w42732;
	assign w42800 = w42819 & w42804;
	assign w42734 = w42800 ^ w42730;
	assign w42797 = w42818 & w42807;
	assign w42733 = w42797 ^ w42731;
	assign w42739 = w42735 ^ w42733;
	assign w42744 = w46405 ^ w42739;
	assign w42705 = w42796 ^ w42797;
	assign w42752 = w42705 ^ w42706;
	assign w42751 = w42752 ^ w42734;
	assign w42795 = w42817 & w42808;
	assign w42894 = w43133 ^ w43129;
	assign w50409 = w50495 ^ w42894;
	assign w46394 = w50409 ^ w410;
	assign w42858 = w43082 ^ w45662;
	assign w43154 = w42858 ^ w42859;
	assign w50400 = w43154 ^ w43140;
	assign w46403 = w50400 ^ w401;
	assign w41791 = w46403 ^ w46401;
	assign w41793 = w46402 ^ w41791;
	assign w41869 = w46398 ^ w41793;
	assign w41866 = w46399 ^ w41793;
	assign w41872 = w41791 ^ w41880;
	assign w41808 = w46403 ^ w46402;
	assign w41876 = w41880 ^ w41808;
	assign w41870 = w41791 ^ w41754;
	assign w41881 = w46397 ^ w46403;
	assign w41865 = w41872 & w41876;
	assign w41797 = w41865 ^ w41794;
	assign w41862 = w41881 & w41866;
	assign w41796 = w41862 ^ w41792;
	assign w41859 = w41880 & w41869;
	assign w41795 = w41859 ^ w41793;
	assign w41801 = w41797 ^ w41795;
	assign w41806 = w46397 ^ w41801;
	assign w41767 = w41858 ^ w41859;
	assign w41814 = w41767 ^ w41768;
	assign w41813 = w41814 ^ w41796;
	assign w41857 = w41879 & w41870;
	assign w39467 = w46389 ^ w46394;
	assign w45663 = ~w29290;
	assign w43137 = w45294 ^ w45663;
	assign w42939 = w43137 ^ w43083;
	assign w50383 = w45763 ^ w42939;
	assign w42924 = w43137 ^ w43078;
	assign w50391 = w45286 ^ w42924;
	assign w50399 = w45663 ^ w42910;
	assign w42898 = w43140 ^ w43137;
	assign w42896 = ~w42898;
	assign w42850 = w42852 ^ w45663;
	assign w43157 = w42850 ^ w42851;
	assign w50384 = w43157 ^ w43129;
	assign w46419 = w50384 ^ w385;
	assign w41925 = w46419 ^ w46417;
	assign w42006 = w41925 ^ w42014;
	assign w42004 = w41925 ^ w41888;
	assign w42015 = w46413 ^ w46419;
	assign w46412 = w50391 ^ w392;
	assign w42809 = w46412 ^ w42810;
	assign w42736 = w46412 ^ w46406;
	assign w42806 = w42736 ^ w42731;
	assign w42813 = w42730 ^ w42736;
	assign w42811 = w42746 ^ w42813;
	assign w42816 = w46407 ^ w42736;
	assign w42812 = w46411 ^ w42816;
	assign w42815 = w46412 ^ w42691;
	assign w42802 = w42811 & w42809;
	assign w42753 = w42796 ^ w42802;
	assign w42794 = w42753 ^ w42744;
	assign w42801 = w46412 & w42815;
	assign w42799 = w42816 & w42812;
	assign w42793 = w42799 ^ w42751;
	assign w42798 = w42813 & w42806;
	assign w42790 = w42794 & w42793;
	assign w46404 = w50399 ^ w400;
	assign w41871 = w46404 ^ w41872;
	assign w41798 = w46404 ^ w46398;
	assign w41868 = w41798 ^ w41793;
	assign w41875 = w41792 ^ w41798;
	assign w41873 = w41808 ^ w41875;
	assign w41878 = w46399 ^ w41798;
	assign w41874 = w46403 ^ w41878;
	assign w41877 = w46404 ^ w41753;
	assign w41864 = w41873 & w41871;
	assign w41815 = w41858 ^ w41864;
	assign w41856 = w41815 ^ w41806;
	assign w41863 = w46404 & w41877;
	assign w41861 = w41878 & w41874;
	assign w41855 = w41861 ^ w41813;
	assign w41860 = w41875 & w41868;
	assign w41852 = w41856 & w41855;
	assign w46420 = w50383 ^ w384;
	assign w42005 = w46420 ^ w42006;
	assign w41932 = w46420 ^ w46414;
	assign w42009 = w41926 ^ w41932;
	assign w42012 = w46415 ^ w41932;
	assign w42008 = w46419 ^ w42012;
	assign w42011 = w46420 ^ w41887;
	assign w41997 = w46420 & w42011;
	assign w41995 = w42012 & w42008;
	assign w45122 = w41857 ^ w41863;
	assign w41807 = w45122 ^ w41792;
	assign w41853 = w41815 ^ w41807;
	assign w41769 = w41801 ^ w45122;
	assign w41812 = w46399 ^ w41769;
	assign w41847 = w41852 ^ w41812;
	assign w45123 = w41857 ^ w41860;
	assign w41810 = w41858 ^ w45123;
	assign w41766 = w41861 ^ w41810;
	assign w41848 = w46403 ^ w41766;
	assign w41846 = w41847 & w41848;
	assign w41844 = w41852 ^ w41846;
	assign w41765 = w41846 ^ w41810;
	assign w41764 = w41846 ^ w41863;
	assign w41759 = w41764 ^ w41860;
	assign w41770 = w41796 ^ w45123;
	assign w41854 = w41770 ^ w41795;
	assign w41845 = w41846 ^ w41854;
	assign w41851 = w41852 ^ w41854;
	assign w41850 = w41853 & w41851;
	assign w41849 = w41850 ^ w41812;
	assign w41761 = w41850 ^ w41862;
	assign w41757 = w41761 ^ w41797;
	assign w41760 = w46397 ^ w41757;
	assign w41837 = w41759 ^ w41760;
	assign w41758 = w41850 ^ w41806;
	assign w41756 = w46399 ^ w41757;
	assign w41843 = w41854 & w41844;
	assign w41841 = w41843 ^ w41851;
	assign w41840 = w41849 & w41841;
	assign w41805 = w41840 ^ w41815;
	assign w41839 = w41805 ^ w41807;
	assign w41763 = w41840 ^ w41864;
	assign w41836 = w41805 ^ w41758;
	assign w41831 = w41845 & w46404;
	assign w41830 = w41836 & w41866;
	assign w41829 = w41839 & w41878;
	assign w41828 = w41849 & w41868;
	assign w41772 = w41828 ^ w41829;
	assign w41827 = w41837 & w41869;
	assign w41822 = w41845 & w41877;
	assign w41821 = w41836 & w41881;
	assign w41788 = w41830 ^ w41821;
	assign w41820 = w41839 & w41874;
	assign w41790 = w41828 ^ w41820;
	assign w41819 = w41849 & w41875;
	assign w41818 = w41837 & w41880;
	assign w45124 = w41829 ^ w41830;
	assign w45126 = w41843 ^ w41861;
	assign w41802 = w46403 ^ w45126;
	assign w41755 = w41802 ^ w41763;
	assign w41762 = w41792 ^ w41755;
	assign w41838 = w41759 ^ w41762;
	assign w41825 = w41838 & w41870;
	assign w41803 = w41821 ^ w41825;
	assign w41781 = ~w41803;
	assign w41834 = w41755 ^ w41756;
	assign w41826 = w41834 & w41867;
	assign w41783 = w41826 ^ w41827;
	assign w41787 = w41826 ^ w41829;
	assign w41784 = ~w41787;
	assign w41780 = w41781 ^ w41819;
	assign w41817 = w41834 & w41882;
	assign w41816 = w41838 & w41879;
	assign w41782 = w41827 ^ w41816;
	assign w41778 = ~w41782;
	assign w43615 = w41817 ^ w41818;
	assign w41786 = w41790 ^ w43615;
	assign w41785 = w41781 ^ w41786;
	assign w41885 = w41784 ^ w41785;
	assign w41842 = w41802 ^ w41765;
	assign w41832 = w41842 & w41871;
	assign w41823 = w41842 & w41873;
	assign w41799 = w41823 ^ w43615;
	assign w41811 = w41826 ^ w45124;
	assign w41777 = w41822 ^ w41811;
	assign w41774 = ~w41777;
	assign w41771 = w41827 ^ w41811;
	assign w41835 = w45126 ^ w41813;
	assign w41833 = w41835 & w41872;
	assign w41824 = w41835 & w41876;
	assign w41800 = w41824 ^ w41799;
	assign w41804 = w41832 ^ w41800;
	assign w41809 = w41833 ^ w41804;
	assign w50715 = w45124 ^ w41809;
	assign w41884 = w41809 ^ w41783;
	assign w41773 = w41831 ^ w41804;
	assign w50714 = w41772 ^ w41773;
	assign w50716 = w41800 ^ w41771;
	assign w9822 = w50716 ^ w50720;
	assign w9798 = w9887 ^ w9822;
	assign w9630 = w50715 ^ w50714;
	assign w9791 = w9857 ^ w50715;
	assign w9842 = w50710 ^ w50714;
	assign w9793 = w9888 ^ w9842;
	assign w50619 = w9910 ^ w9842;
	assign w46257 = w50619 ^ w483;
	assign w9837 = w50712 ^ w50716;
	assign w9794 = w9837 ^ w50719;
	assign w50636 = w9793 ^ w9794;
	assign w46240 = w50636 ^ w500;
	assign w9806 = w45951 ^ w50714;
	assign w50627 = w9805 ^ w9806;
	assign w46249 = w50627 ^ w491;
	assign w9797 = w9885 ^ w9837;
	assign w50632 = w45828 ^ w9797;
	assign w46244 = w50632 ^ w496;
	assign w9574 = w9837 ^ w45827;
	assign w9839 = w50715 ^ w50719;
	assign w9819 = w9848 ^ w9839;
	assign w50620 = w9819 ^ w9820;
	assign w9787 = w9885 ^ w9822;
	assign w45125 = w41831 ^ w41833;
	assign w41789 = w45125 ^ w41786;
	assign w41886 = w41788 ^ w41789;
	assign w41776 = w41780 ^ w45125;
	assign w41779 = w41818 ^ w41776;
	assign w41883 = w41778 ^ w41779;
	assign w41775 = w41799 ^ w41776;
	assign w50713 = w41774 ^ w41775;
	assign w9840 = w50713 ^ w50717;
	assign w9631 = w9840 ^ w45576;
	assign w9576 = w9837 ^ w50713;
	assign w9916 = w9576 ^ w9577;
	assign w50618 = w9631 ^ w9632;
	assign w9808 = w9877 ^ w9840;
	assign w50626 = w50704 ^ w9808;
	assign w46250 = w50626 ^ w490;
	assign w40428 = w46249 ^ w46250;
	assign w45161 = w42795 ^ w42801;
	assign w42745 = w45161 ^ w42730;
	assign w42791 = w42753 ^ w42745;
	assign w42707 = w42739 ^ w45161;
	assign w42750 = w46407 ^ w42707;
	assign w42785 = w42790 ^ w42750;
	assign w45162 = w42795 ^ w42798;
	assign w42748 = w42796 ^ w45162;
	assign w42704 = w42799 ^ w42748;
	assign w42786 = w46411 ^ w42704;
	assign w42784 = w42785 & w42786;
	assign w42703 = w42784 ^ w42748;
	assign w42702 = w42784 ^ w42801;
	assign w42697 = w42702 ^ w42798;
	assign w42782 = w42790 ^ w42784;
	assign w42708 = w42734 ^ w45162;
	assign w42792 = w42708 ^ w42733;
	assign w42783 = w42784 ^ w42792;
	assign w42789 = w42790 ^ w42792;
	assign w42788 = w42789 & w42791;
	assign w42787 = w42788 ^ w42750;
	assign w42699 = w42788 ^ w42800;
	assign w42695 = w42699 ^ w42735;
	assign w42698 = w46405 ^ w42695;
	assign w42775 = w42697 ^ w42698;
	assign w42696 = w42788 ^ w42744;
	assign w42694 = w46407 ^ w42695;
	assign w42781 = w42792 & w42782;
	assign w42779 = w42781 ^ w42789;
	assign w42778 = w42787 & w42779;
	assign w42743 = w42778 ^ w42753;
	assign w42777 = w42743 ^ w42745;
	assign w42701 = w42778 ^ w42802;
	assign w42774 = w42743 ^ w42696;
	assign w42769 = w42783 & w46412;
	assign w42768 = w42774 & w42804;
	assign w42767 = w42777 & w42816;
	assign w42766 = w42787 & w42806;
	assign w42710 = w42766 ^ w42767;
	assign w42765 = w42775 & w42807;
	assign w42760 = w42783 & w42815;
	assign w42759 = w42774 & w42819;
	assign w42726 = w42768 ^ w42759;
	assign w42758 = w42777 & w42812;
	assign w42728 = w42766 ^ w42758;
	assign w42757 = w42787 & w42813;
	assign w42756 = w42775 & w42818;
	assign w45163 = w42767 ^ w42768;
	assign w45165 = w42781 ^ w42799;
	assign w42740 = w46411 ^ w45165;
	assign w42780 = w42740 ^ w42703;
	assign w42761 = w42780 & w42811;
	assign w42770 = w42780 & w42809;
	assign w42693 = w42740 ^ w42701;
	assign w42700 = w42730 ^ w42693;
	assign w42776 = w42697 ^ w42700;
	assign w42763 = w42776 & w42808;
	assign w42741 = w42759 ^ w42763;
	assign w42719 = ~w42741;
	assign w42718 = w42719 ^ w42757;
	assign w42772 = w42693 ^ w42694;
	assign w42755 = w42772 & w42820;
	assign w42754 = w42776 & w42817;
	assign w42720 = w42765 ^ w42754;
	assign w42716 = ~w42720;
	assign w43618 = w42755 ^ w42756;
	assign w42737 = w42761 ^ w43618;
	assign w42724 = w42728 ^ w43618;
	assign w42723 = w42719 ^ w42724;
	assign w42764 = w42772 & w42805;
	assign w42725 = w42764 ^ w42767;
	assign w42722 = ~w42725;
	assign w42823 = w42722 ^ w42723;
	assign w42721 = w42764 ^ w42765;
	assign w42749 = w42764 ^ w45163;
	assign w42709 = w42765 ^ w42749;
	assign w42715 = w42760 ^ w42749;
	assign w42712 = ~w42715;
	assign w42773 = w45165 ^ w42751;
	assign w42771 = w42773 & w42810;
	assign w42762 = w42773 & w42814;
	assign w42738 = w42762 ^ w42737;
	assign w42742 = w42770 ^ w42738;
	assign w42747 = w42771 ^ w42742;
	assign w50654 = w45163 ^ w42747;
	assign w42822 = w42747 ^ w42721;
	assign w42711 = w42769 ^ w42742;
	assign w50653 = w42710 ^ w42711;
	assign w9893 = w50649 ^ w50653;
	assign w50657 = w42738 ^ w42709;
	assign w50656 = ~w42822;
	assign w9731 = w9732 ^ w50653;
	assign w50523 = w9730 ^ w9731;
	assign w9616 = w50660 ^ w50653;
	assign w9758 = w50661 ^ w50654;
	assign w46353 = w50523 ^ w578;
	assign w9884 = w50650 ^ w50654;
	assign w9681 = w45509 ^ w42822;
	assign w9679 = w9680 ^ w9681;
	assign w50547 = w9896 ^ w9893;
	assign w9772 = w9884 ^ w9876;
	assign w50526 = ~w9679;
	assign w46350 = w50526 ^ w581;
	assign w50533 = w45278 ^ w9772;
	assign w46343 = w50533 ^ w588;
	assign w9748 = w9884 ^ w9883;
	assign w9746 = ~w9748;
	assign w50548 = w9746 ^ w9747;
	assign w46329 = w50547 ^ w602;
	assign w46328 = w50548 ^ w603;
	assign w9829 = w50651 ^ w50657;
	assign w9644 = w9892 ^ w9829;
	assign w9619 = w9829 ^ w50649;
	assign w9742 = w9873 ^ w9829;
	assign w50551 = w50662 ^ w9742;
	assign w46325 = w50551 ^ w606;
	assign w39334 = w46328 ^ w46325;
	assign w50528 = w45864 ^ w9644;
	assign w46348 = w50528 ^ w583;
	assign w45164 = w42769 ^ w42771;
	assign w42727 = w45164 ^ w42724;
	assign w42824 = w42726 ^ w42727;
	assign w42714 = w42718 ^ w45164;
	assign w42717 = w42756 ^ w42714;
	assign w42821 = w42716 ^ w42717;
	assign w42713 = w42737 ^ w42714;
	assign w50652 = w42712 ^ w42713;
	assign w50655 = ~w42821;
	assign w9620 = w50648 ^ w50652;
	assign w9868 = w50652 ^ w50659;
	assign w9898 = w9619 ^ w9620;
	assign w9751 = ~w9868;
	assign w9881 = w45278 ^ w50655;
	assign w9771 = w9881 ^ w9873;
	assign w9757 = w9881 ^ w45509;
	assign w50541 = w9757 ^ w9758;
	assign w46335 = w50541 ^ w596;
	assign w9744 = w9891 ^ w9868;
	assign w9762 = w9893 ^ w9751;
	assign w9745 = w9881 ^ w9880;
	assign w50549 = w45862 ^ w9745;
	assign w46327 = w50549 ^ w604;
	assign w39246 = w46327 ^ w46325;
	assign w9698 = w50665 ^ w42821;
	assign w50534 = w45279 ^ w9771;
	assign w50522 = w50663 ^ w9744;
	assign w46354 = w50522 ^ w577;
	assign w41500 = w46353 ^ w46354;
	assign w46342 = w50534 ^ w589;
	assign w40726 = w46348 ^ w46342;
	assign w40806 = w46343 ^ w40726;
	assign w50525 = w9697 ^ w9698;
	assign w46258 = w50618 ^ w482;
	assign w41098 = w46257 ^ w46258;
	assign w50635 = w9916 ^ w9848;
	assign w46241 = w50635 ^ w499;
	assign w9879 = w45279 ^ w50656;
	assign w9743 = w9879 ^ w9876;
	assign w9755 = w9879 ^ w23526;
	assign w9770 = w9879 ^ w9828;
	assign w50550 = w45863 ^ w9743;
	assign w46326 = w50550 ^ w605;
	assign w39248 = w46328 ^ w46326;
	assign w39208 = w39248 ^ w39246;
	assign w39207 = w39248 ^ w46327;
	assign w9775 = ~w9893;
	assign w9773 = w9775 ^ w9880;
	assign w50531 = w9898 ^ w9883;
	assign w50535 = w50651 ^ w9770;
	assign w46341 = w50535 ^ w590;
	assign w40720 = w46343 ^ w46341;
	assign w40803 = w40720 ^ w40726;
	assign w9629 = w9822 ^ w50718;
	assign w9894 = w9629 ^ w9630;
	assign w50644 = w9894 ^ w9888;
	assign w9756 = w45862 ^ w42821;
	assign w50542 = w9755 ^ w9756;
	assign w46334 = w50542 ^ w597;
	assign w50631 = w50708 ^ w9798;
	assign w46245 = w50631 ^ w495;
	assign w40539 = w46245 ^ w46250;
	assign w9749 = w9751 ^ w50648;
	assign w50546 = w9749 ^ w9750;
	assign w46330 = w50546 ^ w601;
	assign w39222 = w46329 ^ w46330;
	assign w39336 = w46330 ^ w46328;
	assign w39321 = w39246 ^ w39336;
	assign w39312 = w39336 & w39321;
	assign w39333 = w46325 ^ w46330;
	assign w9661 = w23526 ^ w50657;
	assign w50527 = w9660 ^ w9661;
	assign w46349 = w50527 ^ w582;
	assign w41611 = w46349 ^ w46354;
	assign w50637 = w9791 ^ w9792;
	assign w46239 = w50637 ^ w501;
	assign w9830 = w50657 ^ w50662;
	assign w9769 = w9892 ^ w9830;
	assign w9615 = w9830 ^ w50665;
	assign w9764 = ~w9830;
	assign w9900 = w9615 ^ w9616;
	assign w9763 = w9764 ^ w50664;
	assign w50539 = w9762 ^ w9763;
	assign w46337 = w50539 ^ w594;
	assign w46351 = w50525 ^ w580;
	assign w41524 = w46351 ^ w46349;
	assign w50628 = w9895 ^ w9839;
	assign w46248 = w50628 ^ w492;
	assign w40540 = w46248 ^ w46245;
	assign w40542 = w46250 ^ w46248;
	assign w46418 = w50385 ^ w386;
	assign w41927 = w46418 ^ w41925;
	assign w42003 = w46414 ^ w41927;
	assign w42000 = w46415 ^ w41927;
	assign w42002 = w41932 ^ w41927;
	assign w41942 = w46419 ^ w46418;
	assign w42007 = w41942 ^ w42009;
	assign w42010 = w42014 ^ w41942;
	assign w42016 = w46418 ^ w46416;
	assign w42001 = w41926 ^ w42016;
	assign w41902 = w46417 ^ w46418;
	assign w42013 = w46413 ^ w46418;
	assign w41999 = w42006 & w42010;
	assign w41931 = w41999 ^ w41928;
	assign w41998 = w42007 & w42005;
	assign w41996 = w42015 & w42000;
	assign w41930 = w41996 ^ w41926;
	assign w41994 = w42009 & w42002;
	assign w41993 = w42014 & w42003;
	assign w41929 = w41993 ^ w41927;
	assign w41935 = w41931 ^ w41929;
	assign w41940 = w46413 ^ w41935;
	assign w41992 = w42016 & w42001;
	assign w41949 = w41992 ^ w41998;
	assign w41990 = w41949 ^ w41940;
	assign w41901 = w41992 ^ w41993;
	assign w41948 = w41901 ^ w41902;
	assign w41947 = w41948 ^ w41930;
	assign w41989 = w41995 ^ w41947;
	assign w41991 = w42013 & w42004;
	assign w41986 = w41990 & w41989;
	assign w45127 = w41991 ^ w41997;
	assign w41903 = w41935 ^ w45127;
	assign w41946 = w46415 ^ w41903;
	assign w41981 = w41986 ^ w41946;
	assign w41941 = w45127 ^ w41926;
	assign w41987 = w41949 ^ w41941;
	assign w45128 = w41991 ^ w41994;
	assign w41944 = w41992 ^ w45128;
	assign w41900 = w41995 ^ w41944;
	assign w41982 = w46419 ^ w41900;
	assign w41980 = w41981 & w41982;
	assign w41899 = w41980 ^ w41944;
	assign w41978 = w41986 ^ w41980;
	assign w41898 = w41980 ^ w41997;
	assign w41893 = w41898 ^ w41994;
	assign w41904 = w41930 ^ w45128;
	assign w41988 = w41904 ^ w41929;
	assign w41979 = w41980 ^ w41988;
	assign w41985 = w41986 ^ w41988;
	assign w41984 = w41987 & w41985;
	assign w41983 = w41984 ^ w41946;
	assign w41895 = w41984 ^ w41996;
	assign w41891 = w41895 ^ w41931;
	assign w41894 = w46413 ^ w41891;
	assign w41971 = w41893 ^ w41894;
	assign w41892 = w41984 ^ w41940;
	assign w41890 = w46415 ^ w41891;
	assign w41977 = w41988 & w41978;
	assign w41975 = w41977 ^ w41985;
	assign w41974 = w41983 & w41975;
	assign w41939 = w41974 ^ w41949;
	assign w41973 = w41939 ^ w41941;
	assign w41897 = w41974 ^ w41998;
	assign w41970 = w41939 ^ w41892;
	assign w41965 = w41979 & w46420;
	assign w41964 = w41970 & w42000;
	assign w41963 = w41973 & w42012;
	assign w41962 = w41983 & w42002;
	assign w41906 = w41962 ^ w41963;
	assign w41961 = w41971 & w42003;
	assign w41956 = w41979 & w42011;
	assign w41955 = w41970 & w42015;
	assign w41922 = w41964 ^ w41955;
	assign w41954 = w41973 & w42008;
	assign w41924 = w41962 ^ w41954;
	assign w41953 = w41983 & w42009;
	assign w41952 = w41971 & w42014;
	assign w45130 = w41963 ^ w41964;
	assign w45132 = w41977 ^ w41995;
	assign w41969 = w45132 ^ w41947;
	assign w41967 = w41969 & w42006;
	assign w45131 = w41965 ^ w41967;
	assign w41958 = w41969 & w42010;
	assign w41936 = w46419 ^ w45132;
	assign w41976 = w41936 ^ w41899;
	assign w41889 = w41936 ^ w41897;
	assign w41896 = w41926 ^ w41889;
	assign w41972 = w41893 ^ w41896;
	assign w41968 = w41889 ^ w41890;
	assign w41966 = w41976 & w42005;
	assign w41960 = w41968 & w42001;
	assign w41945 = w41960 ^ w45130;
	assign w41921 = w41960 ^ w41963;
	assign w41918 = ~w41921;
	assign w41917 = w41960 ^ w41961;
	assign w41911 = w41956 ^ w41945;
	assign w41908 = ~w41911;
	assign w41905 = w41961 ^ w41945;
	assign w41959 = w41972 & w42004;
	assign w41937 = w41955 ^ w41959;
	assign w41915 = ~w41937;
	assign w41914 = w41915 ^ w41953;
	assign w41910 = w41914 ^ w45131;
	assign w41913 = w41952 ^ w41910;
	assign w41957 = w41976 & w42007;
	assign w41951 = w41968 & w42016;
	assign w41950 = w41972 & w42013;
	assign w41916 = w41961 ^ w41950;
	assign w41912 = ~w41916;
	assign w42017 = w41912 ^ w41913;
	assign w45129 = w41951 ^ w41952;
	assign w41933 = w41957 ^ w45129;
	assign w41909 = w41933 ^ w41910;
	assign w50668 = w41908 ^ w41909;
	assign w41934 = w41958 ^ w41933;
	assign w50671 = w41934 ^ w41905;
	assign w41938 = w41966 ^ w41934;
	assign w41907 = w41965 ^ w41938;
	assign w50669 = w41906 ^ w41907;
	assign w9858 = w50669 ^ w50674;
	assign w41943 = w41967 ^ w41938;
	assign w42018 = w41943 ^ w41917;
	assign w50571 = w9908 ^ w9858;
	assign w9587 = w50675 ^ w50669;
	assign w9584 = w9585 ^ w50668;
	assign w9722 = ~w9858;
	assign w9720 = w9722 ^ w9846;
	assign w9861 = w50668 ^ w50673;
	assign w9702 = w9861 ^ w9859;
	assign w9714 = ~w9861;
	assign w9712 = w9714 ^ w50681;
	assign w9826 = w50671 ^ w50676;
	assign w9706 = w9843 ^ w9826;
	assign w50575 = w50684 ^ w9706;
	assign w9700 = w9858 ^ w9856;
	assign w50579 = w9700 ^ w9701;
	assign w46297 = w50579 ^ w570;
	assign w9723 = w9714 ^ w9851;
	assign w50570 = w9712 ^ w9713;
	assign w46306 = w50570 ^ w561;
	assign w9689 = w9826 ^ w45818;
	assign w50583 = w9689 ^ w9690;
	assign w50578 = w50677 ^ w9702;
	assign w46298 = w50578 ^ w569;
	assign w39088 = w46297 ^ w46298;
	assign w50670 = w45130 ^ w41943;
	assign w9854 = w50670 ^ w50675;
	assign w9719 = w9854 ^ w9841;
	assign w9738 = w45848 ^ w50670;
	assign w50557 = w9737 ^ w9738;
	assign w50572 = w9907 ^ w9854;
	assign w46304 = w50572 ^ w563;
	assign w41480 = w46306 ^ w46304;
	assign w46319 = w50557 ^ w548;
	assign w41920 = w41924 ^ w45129;
	assign w41923 = w45131 ^ w41920;
	assign w42020 = w41922 ^ w41923;
	assign w41919 = w41915 ^ w41920;
	assign w42019 = w41918 ^ w41919;
	assign w46301 = w50575 ^ w566;
	assign w41478 = w46304 ^ w46301;
	assign w41477 = w46301 ^ w46306;
	assign w46305 = w50571 ^ w562;
	assign w41366 = w46305 ^ w46306;
	assign w9835 = w50671 ^ w50684;
	assign w9582 = ~w9835;
	assign w9583 = w9582 ^ w50681;
	assign w9913 = w9583 ^ w9584;
	assign w50555 = w9913 ^ w9851;
	assign w46321 = w50555 ^ w546;
	assign w9586 = w9835 ^ w50682;
	assign w9912 = w9586 ^ w9587;
	assign w50556 = w9912 ^ w9846;
	assign w46320 = w50556 ^ w547;
	assign w9741 = w9863 ^ w9835;
	assign w50552 = w45842 ^ w9741;
	assign w46324 = w50552 ^ w543;
	assign w9729 = w9863 ^ w9826;
	assign w9580 = w9582 ^ w45820;
	assign w46293 = w50583 ^ w574;
	assign w39199 = w46293 ^ w46298;
	assign w9696 = ~w9854;
	assign w9693 = w9696 ^ w9851;
	assign w50580 = w9693 ^ w9694;
	assign w46296 = w50580 ^ w571;
	assign w39202 = w46298 ^ w46296;
	assign w39200 = w46296 ^ w46293;
	assign w9781 = w9842 ^ w9840;
	assign w45866 = ~w41883;
	assign w9847 = w45215 ^ w45866;
	assign w9779 = w9847 ^ w9839;
	assign w9818 = ~w9847;
	assign w9816 = w9818 ^ w45833;
	assign w50621 = w9816 ^ w9817;
	assign w46255 = w50621 ^ w485;
	assign w50629 = w45866 ^ w9804;
	assign w46247 = w50629 ^ w493;
	assign w40452 = w46247 ^ w46245;
	assign w40527 = w40452 ^ w40542;
	assign w40518 = w40542 & w40527;
	assign w50645 = w45575 ^ w9779;
	assign w46231 = w50645 ^ w45168;
	assign w9790 = w9887 ^ w9847;
	assign w50638 = w45826 ^ w9790;
	assign w46238 = w50638 ^ w502;
	assign w42330 = w46240 ^ w46238;
	assign w42334 = w46244 ^ w46238;
	assign w42414 = w46239 ^ w42334;
	assign w42289 = w42330 ^ w46239;
	assign w42413 = w46244 ^ w42289;
	assign w42399 = w46244 & w42413;
	assign w45867 = ~w41884;
	assign w9845 = w45867 ^ w45826;
	assign w9800 = w9845 ^ w45215;
	assign w9815 = w9857 ^ w9845;
	assign w50622 = w45216 ^ w9815;
	assign w46254 = w50622 ^ w486;
	assign w9789 = w45867 ^ w45216;
	assign w50639 = w9788 ^ w9789;
	assign w46237 = w50639 ^ w503;
	assign w42328 = w46239 ^ w46237;
	assign w42416 = w46240 ^ w46237;
	assign w42411 = w42328 ^ w42334;
	assign w42290 = w42330 ^ w42328;
	assign w9778 = w45867 ^ w45866;
	assign w50646 = w9777 ^ w9778;
	assign w9776 = w9845 ^ w9823;
	assign w50647 = w50716 ^ w9776;
	assign w46229 = w50647 ^ w510;
	assign w38978 = w46231 ^ w46229;
	assign w46230 = w50646 ^ w509;
	assign w9799 = w9800 ^ w9801;
	assign w50630 = ~w9799;
	assign w46246 = w50630 ^ w494;
	assign w40454 = w46248 ^ w46246;
	assign w40414 = w40454 ^ w40452;
	assign w40413 = w40454 ^ w46247;
	assign w45868 = ~w41885;
	assign w9852 = w45868 ^ w45827;
	assign w9783 = w9862 ^ w9852;
	assign w50617 = w9911 ^ w9852;
	assign w46259 = w50617 ^ w481;
	assign w41121 = w46259 ^ w46257;
	assign w41123 = w46258 ^ w41121;
	assign w41199 = w46254 ^ w41123;
	assign w41196 = w46255 ^ w41123;
	assign w41138 = w46259 ^ w46258;
	assign w9810 = w9885 ^ w9852;
	assign w9809 = w9810 ^ w9811;
	assign w50625 = ~w9809;
	assign w46251 = w50625 ^ w489;
	assign w40451 = w46251 ^ w46249;
	assign w40453 = w46250 ^ w40451;
	assign w40529 = w46246 ^ w40453;
	assign w40526 = w46247 ^ w40453;
	assign w40532 = w40451 ^ w40540;
	assign w40468 = w46251 ^ w46250;
	assign w40536 = w40540 ^ w40468;
	assign w40530 = w40451 ^ w40414;
	assign w40541 = w46245 ^ w46251;
	assign w40525 = w40532 & w40536;
	assign w40457 = w40525 ^ w40454;
	assign w40522 = w40541 & w40526;
	assign w40456 = w40522 ^ w40452;
	assign w40519 = w40540 & w40529;
	assign w40455 = w40519 ^ w40453;
	assign w40461 = w40457 ^ w40455;
	assign w40466 = w46245 ^ w40461;
	assign w40427 = w40518 ^ w40519;
	assign w40474 = w40427 ^ w40428;
	assign w40473 = w40474 ^ w40456;
	assign w40517 = w40539 & w40530;
	assign w50642 = w50713 ^ w9783;
	assign w46234 = w50642 ^ w506;
	assign w39065 = w46229 ^ w46234;
	assign w9796 = w45868 ^ w45217;
	assign w50634 = w9795 ^ w9796;
	assign w46242 = w50634 ^ w498;
	assign w42418 = w46242 ^ w46240;
	assign w42403 = w42328 ^ w42418;
	assign w42304 = w46241 ^ w46242;
	assign w42415 = w46237 ^ w46242;
	assign w42394 = w42418 & w42403;
	assign w45869 = ~w41886;
	assign w50640 = w45869 ^ w9787;
	assign w46236 = w50640 ^ w504;
	assign w38984 = w46236 ^ w46230;
	assign w39061 = w38978 ^ w38984;
	assign w39064 = w46231 ^ w38984;
	assign w9575 = w45869 ^ w45213;
	assign w9917 = w9574 ^ w9575;
	assign w50633 = w9917 ^ w9877;
	assign w46243 = w50633 ^ w497;
	assign w42327 = w46243 ^ w46241;
	assign w42329 = w46242 ^ w42327;
	assign w42405 = w46238 ^ w42329;
	assign w42402 = w46239 ^ w42329;
	assign w42404 = w42334 ^ w42329;
	assign w42410 = w46243 ^ w42414;
	assign w42408 = w42327 ^ w42416;
	assign w42407 = w46244 ^ w42408;
	assign w42344 = w46243 ^ w46242;
	assign w42409 = w42344 ^ w42411;
	assign w42412 = w42416 ^ w42344;
	assign w42406 = w42327 ^ w42290;
	assign w42417 = w46237 ^ w46243;
	assign w42401 = w42408 & w42412;
	assign w42333 = w42401 ^ w42330;
	assign w42400 = w42409 & w42407;
	assign w42351 = w42394 ^ w42400;
	assign w42398 = w42417 & w42402;
	assign w42332 = w42398 ^ w42328;
	assign w42397 = w42414 & w42410;
	assign w42396 = w42411 & w42404;
	assign w42395 = w42416 & w42405;
	assign w42331 = w42395 ^ w42329;
	assign w42337 = w42333 ^ w42331;
	assign w42342 = w46237 ^ w42337;
	assign w42392 = w42351 ^ w42342;
	assign w42303 = w42394 ^ w42395;
	assign w42350 = w42303 ^ w42304;
	assign w42349 = w42350 ^ w42332;
	assign w42391 = w42397 ^ w42349;
	assign w42393 = w42415 & w42406;
	assign w42388 = w42392 & w42391;
	assign w45144 = w42393 ^ w42399;
	assign w42305 = w42337 ^ w45144;
	assign w42348 = w46239 ^ w42305;
	assign w42383 = w42388 ^ w42348;
	assign w42343 = w45144 ^ w42328;
	assign w42389 = w42351 ^ w42343;
	assign w45145 = w42393 ^ w42396;
	assign w42346 = w42394 ^ w45145;
	assign w42302 = w42397 ^ w42346;
	assign w42384 = w46243 ^ w42302;
	assign w42382 = w42383 & w42384;
	assign w42301 = w42382 ^ w42346;
	assign w42380 = w42388 ^ w42382;
	assign w42300 = w42382 ^ w42399;
	assign w42295 = w42300 ^ w42396;
	assign w42306 = w42332 ^ w45145;
	assign w42390 = w42306 ^ w42331;
	assign w42381 = w42382 ^ w42390;
	assign w42387 = w42388 ^ w42390;
	assign w42386 = w42389 & w42387;
	assign w42385 = w42386 ^ w42348;
	assign w42297 = w42386 ^ w42398;
	assign w42293 = w42297 ^ w42333;
	assign w42296 = w46237 ^ w42293;
	assign w42373 = w42295 ^ w42296;
	assign w42294 = w42386 ^ w42342;
	assign w42292 = w46239 ^ w42293;
	assign w42379 = w42390 & w42380;
	assign w42377 = w42379 ^ w42387;
	assign w42376 = w42385 & w42377;
	assign w42341 = w42376 ^ w42351;
	assign w42375 = w42341 ^ w42343;
	assign w42299 = w42376 ^ w42400;
	assign w42372 = w42341 ^ w42294;
	assign w42367 = w42381 & w46244;
	assign w42366 = w42372 & w42402;
	assign w42365 = w42375 & w42414;
	assign w42364 = w42385 & w42404;
	assign w42308 = w42364 ^ w42365;
	assign w42363 = w42373 & w42405;
	assign w42358 = w42381 & w42413;
	assign w42357 = w42372 & w42417;
	assign w42324 = w42366 ^ w42357;
	assign w42356 = w42375 & w42410;
	assign w42326 = w42364 ^ w42356;
	assign w42355 = w42385 & w42411;
	assign w42354 = w42373 & w42416;
	assign w45147 = w42365 ^ w42366;
	assign w45149 = w42379 ^ w42397;
	assign w42371 = w45149 ^ w42349;
	assign w42369 = w42371 & w42408;
	assign w45148 = w42367 ^ w42369;
	assign w42360 = w42371 & w42412;
	assign w42338 = w46243 ^ w45149;
	assign w42378 = w42338 ^ w42301;
	assign w42291 = w42338 ^ w42299;
	assign w42298 = w42328 ^ w42291;
	assign w42374 = w42295 ^ w42298;
	assign w42370 = w42291 ^ w42292;
	assign w42368 = w42378 & w42407;
	assign w42362 = w42370 & w42403;
	assign w42347 = w42362 ^ w45147;
	assign w42323 = w42362 ^ w42365;
	assign w42320 = ~w42323;
	assign w42319 = w42362 ^ w42363;
	assign w42313 = w42358 ^ w42347;
	assign w42310 = ~w42313;
	assign w42307 = w42363 ^ w42347;
	assign w42361 = w42374 & w42406;
	assign w42339 = w42357 ^ w42361;
	assign w42317 = ~w42339;
	assign w42316 = w42317 ^ w42355;
	assign w42312 = w42316 ^ w45148;
	assign w42315 = w42354 ^ w42312;
	assign w42359 = w42378 & w42409;
	assign w42353 = w42370 & w42418;
	assign w42352 = w42374 & w42415;
	assign w42318 = w42363 ^ w42352;
	assign w42314 = ~w42318;
	assign w42419 = w42314 ^ w42315;
	assign w45146 = w42353 ^ w42354;
	assign w42335 = w42359 ^ w45146;
	assign w42311 = w42335 ^ w42312;
	assign w50860 = w42310 ^ w42311;
	assign w42336 = w42360 ^ w42335;
	assign w50863 = w42336 ^ w42307;
	assign w42340 = w42368 ^ w42336;
	assign w42309 = w42367 ^ w42340;
	assign w50861 = w42308 ^ w42309;
	assign w42345 = w42369 ^ w42340;
	assign w42420 = w42345 ^ w42319;
	assign w10238 = ~w50860;
	assign w10237 = w50861 ^ w10238;
	assign w50862 = w45147 ^ w42345;
	assign w42322 = w42326 ^ w45146;
	assign w42325 = w45148 ^ w42322;
	assign w42422 = w42324 ^ w42325;
	assign w42321 = w42317 ^ w42322;
	assign w42421 = w42320 ^ w42321;
	assign w50859 = ~w42421;
	assign w45870 = ~w42017;
	assign w9736 = w45825 ^ w45870;
	assign w50558 = w9735 ^ w9736;
	assign w46318 = w50558 ^ w549;
	assign w9964 = w46324 ^ w46318;
	assign w50565 = w45870 ^ w9719;
	assign w46311 = w50565 ^ w556;
	assign w10044 = w46319 ^ w9964;
	assign w9960 = w46320 ^ w46318;
	assign w9919 = w9960 ^ w46319;
	assign w10043 = w46324 ^ w9919;
	assign w10029 = w46324 & w10043;
	assign w9850 = w45870 ^ w45848;
	assign w9692 = w9850 ^ w9846;
	assign w50581 = w45282 ^ w9692;
	assign w9711 = w9850 ^ w45825;
	assign w9709 = ~w9711;
	assign w50573 = w9709 ^ w9710;
	assign w46303 = w50573 ^ w564;
	assign w41390 = w46303 ^ w46301;
	assign w41465 = w41390 ^ w41480;
	assign w41456 = w41480 & w41465;
	assign w46295 = w50581 ^ w572;
	assign w39112 = w46295 ^ w46293;
	assign w39187 = w39112 ^ w39202;
	assign w39178 = w39202 & w39187;
	assign w45871 = ~w42018;
	assign w9717 = w50671 ^ w45871;
	assign w50582 = w45871 ^ w9691;
	assign w46294 = w50582 ^ w573;
	assign w39114 = w46296 ^ w46294;
	assign w39074 = w39114 ^ w39112;
	assign w39073 = w39114 ^ w46295;
	assign w50567 = w9716 ^ w9717;
	assign w9844 = w45871 ^ w45818;
	assign w9718 = w9850 ^ w9844;
	assign w50566 = w45283 ^ w9718;
	assign w9707 = w9844 ^ w45282;
	assign w46310 = w50566 ^ w557;
	assign w9734 = w9844 ^ w9825;
	assign w50559 = w50676 ^ w9734;
	assign w46317 = w50559 ^ w550;
	assign w10046 = w46320 ^ w46317;
	assign w9958 = w46319 ^ w46317;
	assign w9920 = w9960 ^ w9958;
	assign w10041 = w9958 ^ w9964;
	assign w50574 = w9707 ^ w9708;
	assign w46302 = w50574 ^ w565;
	assign w41392 = w46304 ^ w46302;
	assign w41352 = w41392 ^ w41390;
	assign w41351 = w41392 ^ w46303;
	assign w46309 = w50567 ^ w558;
	assign w10092 = w46311 ^ w46309;
	assign w45872 = ~w42019;
	assign w9865 = w45872 ^ w50672;
	assign w9725 = w9865 ^ w9856;
	assign w50562 = w50668 ^ w9725;
	assign w46314 = w50562 ^ w553;
	assign w10179 = w46309 ^ w46314;
	assign w50569 = w9909 ^ w9865;
	assign w46307 = w50569 ^ w560;
	assign w41389 = w46307 ^ w46305;
	assign w41391 = w46306 ^ w41389;
	assign w41467 = w46302 ^ w41391;
	assign w41464 = w46303 ^ w41391;
	assign w41470 = w41389 ^ w41478;
	assign w41406 = w46307 ^ w46306;
	assign w41474 = w41478 ^ w41406;
	assign w41468 = w41389 ^ w41352;
	assign w41479 = w46301 ^ w46307;
	assign w41463 = w41470 & w41474;
	assign w41395 = w41463 ^ w41392;
	assign w41460 = w41479 & w41464;
	assign w41394 = w41460 ^ w41390;
	assign w41457 = w41478 & w41467;
	assign w41393 = w41457 ^ w41391;
	assign w41399 = w41395 ^ w41393;
	assign w41404 = w46301 ^ w41399;
	assign w41365 = w41456 ^ w41457;
	assign w41412 = w41365 ^ w41366;
	assign w41411 = w41412 ^ w41394;
	assign w41455 = w41477 & w41468;
	assign w9740 = w50673 ^ w45872;
	assign w50554 = w9739 ^ w9740;
	assign w9703 = w9865 ^ w9863;
	assign w50577 = w9703 ^ w9704;
	assign w46299 = w50577 ^ w568;
	assign w39201 = w46293 ^ w46299;
	assign w39111 = w46299 ^ w46297;
	assign w39190 = w39111 ^ w39074;
	assign w39177 = w39199 & w39190;
	assign w39113 = w46298 ^ w39111;
	assign w39189 = w46294 ^ w39113;
	assign w39179 = w39200 & w39189;
	assign w39087 = w39178 ^ w39179;
	assign w39134 = w39087 ^ w39088;
	assign w39115 = w39179 ^ w39113;
	assign w39192 = w39111 ^ w39200;
	assign w39186 = w46295 ^ w39113;
	assign w39182 = w39201 & w39186;
	assign w39116 = w39182 ^ w39112;
	assign w39128 = w46299 ^ w46298;
	assign w39196 = w39200 ^ w39128;
	assign w39185 = w39192 & w39196;
	assign w39133 = w39134 ^ w39116;
	assign w39117 = w39185 ^ w39114;
	assign w39121 = w39117 ^ w39115;
	assign w39126 = w46293 ^ w39121;
	assign w45873 = ~w42020;
	assign w9866 = w45873 ^ w45842;
	assign w9705 = w9866 ^ w9825;
	assign w9715 = w9866 ^ w9833;
	assign w50576 = w45285 ^ w9705;
	assign w9727 = w9866 ^ w9859;
	assign w9581 = w40947 ^ w45873;
	assign w9914 = w9580 ^ w9581;
	assign w50553 = w9914 ^ w9859;
	assign w46323 = w50553 ^ w544;
	assign w10047 = w46317 ^ w46323;
	assign w9957 = w46323 ^ w46321;
	assign w10036 = w9957 ^ w9920;
	assign w10038 = w9957 ^ w10046;
	assign w10037 = w46324 ^ w10038;
	assign w50560 = w45873 ^ w9729;
	assign w46316 = w50560 ^ w551;
	assign w10098 = w46316 ^ w46310;
	assign w10178 = w46311 ^ w10098;
	assign w10175 = w10092 ^ w10098;
	assign w50568 = w45820 ^ w9715;
	assign w46308 = w50568 ^ w559;
	assign w41469 = w46308 ^ w41470;
	assign w41396 = w46308 ^ w46302;
	assign w41466 = w41396 ^ w41391;
	assign w41473 = w41390 ^ w41396;
	assign w41471 = w41406 ^ w41473;
	assign w41476 = w46303 ^ w41396;
	assign w41472 = w46307 ^ w41476;
	assign w41475 = w46308 ^ w41351;
	assign w41462 = w41471 & w41469;
	assign w41413 = w41456 ^ w41462;
	assign w41454 = w41413 ^ w41404;
	assign w41461 = w46308 & w41475;
	assign w41459 = w41476 & w41472;
	assign w41453 = w41459 ^ w41411;
	assign w41458 = w41473 & w41466;
	assign w41450 = w41454 & w41453;
	assign w45106 = w41455 ^ w41461;
	assign w41405 = w45106 ^ w41390;
	assign w41451 = w41413 ^ w41405;
	assign w41367 = w41399 ^ w45106;
	assign w41410 = w46303 ^ w41367;
	assign w41445 = w41450 ^ w41410;
	assign w45107 = w41455 ^ w41458;
	assign w41408 = w41456 ^ w45107;
	assign w41364 = w41459 ^ w41408;
	assign w41446 = w46307 ^ w41364;
	assign w41444 = w41445 & w41446;
	assign w41363 = w41444 ^ w41408;
	assign w41362 = w41444 ^ w41461;
	assign w41357 = w41362 ^ w41458;
	assign w41442 = w41450 ^ w41444;
	assign w41368 = w41394 ^ w45107;
	assign w41452 = w41368 ^ w41393;
	assign w41443 = w41444 ^ w41452;
	assign w41449 = w41450 ^ w41452;
	assign w41448 = w41451 & w41449;
	assign w41447 = w41448 ^ w41410;
	assign w41359 = w41448 ^ w41460;
	assign w41355 = w41359 ^ w41395;
	assign w41358 = w46301 ^ w41355;
	assign w41435 = w41357 ^ w41358;
	assign w41356 = w41448 ^ w41404;
	assign w41354 = w46303 ^ w41355;
	assign w41441 = w41452 & w41442;
	assign w41439 = w41441 ^ w41449;
	assign w41438 = w41447 & w41439;
	assign w41403 = w41438 ^ w41413;
	assign w41437 = w41403 ^ w41405;
	assign w41361 = w41438 ^ w41462;
	assign w41434 = w41403 ^ w41356;
	assign w41429 = w41443 & w46308;
	assign w41428 = w41434 & w41464;
	assign w41427 = w41437 & w41476;
	assign w41426 = w41447 & w41466;
	assign w41370 = w41426 ^ w41427;
	assign w41425 = w41435 & w41467;
	assign w41420 = w41443 & w41475;
	assign w41419 = w41434 & w41479;
	assign w41386 = w41428 ^ w41419;
	assign w41418 = w41437 & w41472;
	assign w41388 = w41426 ^ w41418;
	assign w41417 = w41447 & w41473;
	assign w41416 = w41435 & w41478;
	assign w45108 = w41427 ^ w41428;
	assign w45110 = w41441 ^ w41459;
	assign w41400 = w46307 ^ w45110;
	assign w41440 = w41400 ^ w41363;
	assign w41421 = w41440 & w41471;
	assign w41430 = w41440 & w41469;
	assign w41353 = w41400 ^ w41361;
	assign w41360 = w41390 ^ w41353;
	assign w41436 = w41357 ^ w41360;
	assign w41423 = w41436 & w41468;
	assign w41401 = w41419 ^ w41423;
	assign w41379 = ~w41401;
	assign w41378 = w41379 ^ w41417;
	assign w41432 = w41353 ^ w41354;
	assign w41415 = w41432 & w41480;
	assign w41414 = w41436 & w41477;
	assign w41380 = w41425 ^ w41414;
	assign w41376 = ~w41380;
	assign w43613 = w41415 ^ w41416;
	assign w41384 = w41388 ^ w43613;
	assign w41383 = w41379 ^ w41384;
	assign w41397 = w41421 ^ w43613;
	assign w41424 = w41432 & w41465;
	assign w41381 = w41424 ^ w41425;
	assign w41385 = w41424 ^ w41427;
	assign w41382 = ~w41385;
	assign w41483 = w41382 ^ w41383;
	assign w41409 = w41424 ^ w45108;
	assign w41375 = w41420 ^ w41409;
	assign w41369 = w41425 ^ w41409;
	assign w41372 = ~w41375;
	assign w41433 = w45110 ^ w41411;
	assign w41431 = w41433 & w41470;
	assign w41422 = w41433 & w41474;
	assign w41398 = w41422 ^ w41397;
	assign w41402 = w41430 ^ w41398;
	assign w41407 = w41431 ^ w41402;
	assign w50899 = w45108 ^ w41407;
	assign w41482 = w41407 ^ w41381;
	assign w41371 = w41429 ^ w41402;
	assign w50898 = w41370 ^ w41371;
	assign w50900 = w41398 ^ w41369;
	assign w45109 = w41429 ^ w41431;
	assign w41387 = w45109 ^ w41384;
	assign w41484 = w41386 ^ w41387;
	assign w41374 = w41378 ^ w45109;
	assign w41377 = w41416 ^ w41374;
	assign w41481 = w41376 ^ w41377;
	assign w41373 = w41397 ^ w41374;
	assign w50897 = w41372 ^ w41373;
	assign w46300 = w50576 ^ w567;
	assign w39197 = w46300 ^ w39073;
	assign w39183 = w46300 & w39197;
	assign w39191 = w46300 ^ w39192;
	assign w45010 = w39177 ^ w39183;
	assign w39127 = w45010 ^ w39112;
	assign w39089 = w39121 ^ w45010;
	assign w39132 = w46295 ^ w39089;
	assign w39118 = w46300 ^ w46294;
	assign w39198 = w46295 ^ w39118;
	assign w39195 = w39112 ^ w39118;
	assign w39193 = w39128 ^ w39195;
	assign w39184 = w39193 & w39191;
	assign w39135 = w39178 ^ w39184;
	assign w39188 = w39118 ^ w39113;
	assign w39180 = w39195 & w39188;
	assign w45011 = w39177 ^ w39180;
	assign w39130 = w39178 ^ w45011;
	assign w39090 = w39116 ^ w45011;
	assign w39194 = w46299 ^ w39198;
	assign w39181 = w39198 & w39194;
	assign w39086 = w39181 ^ w39130;
	assign w39168 = w46299 ^ w39086;
	assign w39174 = w39090 ^ w39115;
	assign w39176 = w39135 ^ w39126;
	assign w39175 = w39181 ^ w39133;
	assign w39172 = w39176 & w39175;
	assign w39171 = w39172 ^ w39174;
	assign w39167 = w39172 ^ w39132;
	assign w39166 = w39167 & w39168;
	assign w39085 = w39166 ^ w39130;
	assign w39084 = w39166 ^ w39183;
	assign w39079 = w39084 ^ w39180;
	assign w39164 = w39172 ^ w39166;
	assign w39163 = w39174 & w39164;
	assign w39165 = w39166 ^ w39174;
	assign w39142 = w39165 & w39197;
	assign w39151 = w39165 & w46300;
	assign w39161 = w39163 ^ w39171;
	assign w45014 = w39163 ^ w39181;
	assign w39122 = w46299 ^ w45014;
	assign w39162 = w39122 ^ w39085;
	assign w39143 = w39162 & w39193;
	assign w39152 = w39162 & w39191;
	assign w39155 = w45014 ^ w39133;
	assign w39144 = w39155 & w39196;
	assign w39153 = w39155 & w39192;
	assign w45013 = w39151 ^ w39153;
	assign w39173 = w39135 ^ w39127;
	assign w39170 = w39173 & w39171;
	assign w39081 = w39170 ^ w39182;
	assign w39078 = w39170 ^ w39126;
	assign w39077 = w39081 ^ w39117;
	assign w39080 = w46293 ^ w39077;
	assign w39157 = w39079 ^ w39080;
	assign w39147 = w39157 & w39189;
	assign w39138 = w39157 & w39200;
	assign w39076 = w46295 ^ w39077;
	assign w39169 = w39170 ^ w39132;
	assign w39139 = w39169 & w39195;
	assign w39160 = w39169 & w39161;
	assign w39125 = w39160 ^ w39135;
	assign w39156 = w39125 ^ w39078;
	assign w39141 = w39156 & w39201;
	assign w39083 = w39160 ^ w39184;
	assign w39150 = w39156 & w39186;
	assign w39075 = w39122 ^ w39083;
	assign w39082 = w39112 ^ w39075;
	assign w39158 = w39079 ^ w39082;
	assign w39145 = w39158 & w39190;
	assign w39123 = w39141 ^ w39145;
	assign w39136 = w39158 & w39199;
	assign w39154 = w39075 ^ w39076;
	assign w39146 = w39154 & w39187;
	assign w39137 = w39154 & w39202;
	assign w39148 = w39169 & w39188;
	assign w39159 = w39125 ^ w39127;
	assign w39149 = w39159 & w39198;
	assign w39140 = w39159 & w39194;
	assign w39110 = w39148 ^ w39140;
	assign w39101 = ~w39123;
	assign w39103 = w39146 ^ w39147;
	assign w39102 = w39147 ^ w39136;
	assign w39098 = ~w39102;
	assign w39108 = w39150 ^ w39141;
	assign w39092 = w39148 ^ w39149;
	assign w43607 = w39137 ^ w39138;
	assign w39119 = w39143 ^ w43607;
	assign w39106 = w39110 ^ w43607;
	assign w39109 = w45013 ^ w39106;
	assign w39100 = w39101 ^ w39139;
	assign w39096 = w39100 ^ w45013;
	assign w39095 = w39119 ^ w39096;
	assign w39099 = w39138 ^ w39096;
	assign w39203 = w39098 ^ w39099;
	assign w45012 = w39149 ^ w39150;
	assign w39131 = w39146 ^ w45012;
	assign w39097 = w39142 ^ w39131;
	assign w39094 = ~w39097;
	assign w50882 = w39094 ^ w39095;
	assign w39091 = w39147 ^ w39131;
	assign w39107 = w39146 ^ w39149;
	assign w39104 = ~w39107;
	assign w39206 = w39108 ^ w39109;
	assign w39105 = w39101 ^ w39106;
	assign w39205 = w39104 ^ w39105;
	assign w39120 = w39144 ^ w39119;
	assign w50885 = w39120 ^ w39091;
	assign w39124 = w39152 ^ w39120;
	assign w39129 = w39153 ^ w39124;
	assign w39093 = w39151 ^ w39124;
	assign w39204 = w39129 ^ w39103;
	assign w50884 = w45012 ^ w39129;
	assign w50883 = w39092 ^ w39093;
	assign w45806 = ~w39205;
	assign w45807 = ~w39206;
	assign w45812 = ~w39203;
	assign w45813 = ~w39204;
	assign w45854 = ~w41483;
	assign w45855 = ~w41484;
	assign w45860 = ~w41481;
	assign w45861 = ~w41482;
	assign w45875 = ~w42419;
	assign w45876 = ~w42420;
	assign w45877 = ~w42422;
	assign w45882 = ~w42824;
	assign w9869 = w45882 ^ w45864;
	assign w9767 = w9891 ^ w9869;
	assign w9752 = w9869 ^ w9828;
	assign w50544 = w45281 ^ w9752;
	assign w9821 = w9869 ^ w9836;
	assign w50520 = w45503 ^ w9821;
	assign w46356 = w50520 ^ w575;
	assign w41530 = w46356 ^ w46350;
	assign w41607 = w41524 ^ w41530;
	assign w41610 = w46351 ^ w41530;
	assign w50536 = w45882 ^ w9769;
	assign w46340 = w50536 ^ w591;
	assign w42602 = w46340 ^ w46334;
	assign w42682 = w46335 ^ w42602;
	assign w46332 = w50544 ^ w599;
	assign w39331 = w46332 ^ w39207;
	assign w39252 = w46332 ^ w46326;
	assign w39332 = w46327 ^ w39252;
	assign w39317 = w46332 & w39331;
	assign w39329 = w39246 ^ w39252;
	assign w45886 = ~w42823;
	assign w9870 = w45886 ^ w50658;
	assign w9802 = w9733 ^ w45886;
	assign w50545 = w9897 ^ w9870;
	assign w46331 = w50545 ^ w600;
	assign w39335 = w46325 ^ w46331;
	assign w39328 = w46331 ^ w39332;
	assign w39245 = w46331 ^ w46329;
	assign w39324 = w39245 ^ w39208;
	assign w39311 = w39333 & w39324;
	assign w39315 = w39332 & w39328;
	assign w50530 = w9802 ^ w9803;
	assign w39262 = w46331 ^ w46330;
	assign w39327 = w39262 ^ w39329;
	assign w39330 = w39334 ^ w39262;
	assign w39247 = w46330 ^ w39245;
	assign w39320 = w46327 ^ w39247;
	assign w39316 = w39335 & w39320;
	assign w39322 = w39252 ^ w39247;
	assign w39323 = w46326 ^ w39247;
	assign w39313 = w39334 & w39323;
	assign w9768 = w9764 ^ w45886;
	assign w9766 = w9767 ^ w9768;
	assign w39249 = w39313 ^ w39247;
	assign w45015 = w39311 ^ w39317;
	assign w39261 = w45015 ^ w39246;
	assign w39250 = w39316 ^ w39246;
	assign w39314 = w39329 & w39322;
	assign w45016 = w39311 ^ w39314;
	assign w39224 = w39250 ^ w45016;
	assign w39308 = w39224 ^ w39249;
	assign w46346 = w50530 ^ w585;
	assign w40807 = w46341 ^ w46346;
	assign w9760 = w9892 ^ w9870;
	assign w9759 = w9760 ^ w9761;
	assign w50521 = ~w9759;
	assign w46355 = w50521 ^ w576;
	assign w41523 = w46355 ^ w46353;
	assign w41525 = w46354 ^ w41523;
	assign w41601 = w46350 ^ w41525;
	assign w41598 = w46351 ^ w41525;
	assign w41600 = w41530 ^ w41525;
	assign w41606 = w46355 ^ w41610;
	assign w41540 = w46355 ^ w46354;
	assign w41605 = w41540 ^ w41607;
	assign w41613 = w46349 ^ w46355;
	assign w41594 = w41613 & w41598;
	assign w41528 = w41594 ^ w41524;
	assign w41593 = w41610 & w41606;
	assign w41592 = w41607 & w41600;
	assign w9765 = w9871 ^ w9870;
	assign w50538 = w50652 ^ w9765;
	assign w46338 = w50538 ^ w593;
	assign w42572 = w46337 ^ w46338;
	assign w50537 = ~w9766;
	assign w46339 = w50537 ^ w592;
	assign w42595 = w46339 ^ w46337;
	assign w42597 = w46338 ^ w42595;
	assign w42673 = w46334 ^ w42597;
	assign w42670 = w46335 ^ w42597;
	assign w42672 = w42602 ^ w42597;
	assign w42678 = w46339 ^ w42682;
	assign w42612 = w46339 ^ w46338;
	assign w42665 = w42682 & w42678;
	assign w39326 = w39245 ^ w39334;
	assign w39325 = w46332 ^ w39326;
	assign w39319 = w39326 & w39330;
	assign w39251 = w39319 ^ w39248;
	assign w39318 = w39327 & w39325;
	assign w39269 = w39312 ^ w39318;
	assign w39307 = w39269 ^ w39261;
	assign w39255 = w39251 ^ w39249;
	assign w39223 = w39255 ^ w45015;
	assign w39266 = w46327 ^ w39223;
	assign w39260 = w46325 ^ w39255;
	assign w39310 = w39269 ^ w39260;
	assign w39264 = w39312 ^ w45016;
	assign w39220 = w39315 ^ w39264;
	assign w39302 = w46331 ^ w39220;
	assign w10040 = w46323 ^ w10044;
	assign w10027 = w10044 & w10040;
	assign w46232 = w50644 ^ w508;
	assign w38980 = w46232 ^ w46230;
	assign w39066 = w46232 ^ w46229;
	assign w39068 = w46234 ^ w46232;
	assign w39053 = w38978 ^ w39068;
	assign w39044 = w39068 & w39053;
	assign w38940 = w38980 ^ w38978;
	assign w38939 = w38980 ^ w46231;
	assign w39063 = w46236 ^ w38939;
	assign w39049 = w46236 & w39063;
	assign w46256 = w50620 ^ w484;
	assign w41124 = w46256 ^ w46254;
	assign w41212 = w46258 ^ w46256;
	assign w41083 = w41124 ^ w46255;
	assign w46345 = w50531 ^ w586;
	assign w40696 = w46345 ^ w46346;
	assign w9872 = w45869 ^ w45828;
	assign w9633 = w9872 ^ w9834;
	assign w9784 = w9786 ^ w9872;
	assign w9812 = w9872 ^ w9823;
	assign w50624 = w45577 ^ w9812;
	assign w46252 = w50624 ^ w488;
	assign w40531 = w46252 ^ w40532;
	assign w40537 = w46252 ^ w40413;
	assign w40523 = w46252 & w40537;
	assign w40458 = w46252 ^ w46246;
	assign w40535 = w40452 ^ w40458;
	assign w40533 = w40468 ^ w40535;
	assign w40524 = w40533 & w40531;
	assign w40475 = w40518 ^ w40524;
	assign w40516 = w40475 ^ w40466;
	assign w40538 = w46247 ^ w40458;
	assign w40534 = w46251 ^ w40538;
	assign w40528 = w40458 ^ w40453;
	assign w40520 = w40535 & w40528;
	assign w40521 = w40538 & w40534;
	assign w40515 = w40521 ^ w40473;
	assign w40512 = w40516 & w40515;
	assign w45066 = w40517 ^ w40523;
	assign w40429 = w40461 ^ w45066;
	assign w40472 = w46247 ^ w40429;
	assign w40507 = w40512 ^ w40472;
	assign w40467 = w45066 ^ w40452;
	assign w40513 = w40475 ^ w40467;
	assign w45067 = w40517 ^ w40520;
	assign w40470 = w40518 ^ w45067;
	assign w40426 = w40521 ^ w40470;
	assign w40508 = w46251 ^ w40426;
	assign w40506 = w40507 & w40508;
	assign w40504 = w40512 ^ w40506;
	assign w40425 = w40506 ^ w40470;
	assign w40424 = w40506 ^ w40523;
	assign w40419 = w40424 ^ w40520;
	assign w40430 = w40456 ^ w45067;
	assign w40514 = w40430 ^ w40455;
	assign w40503 = w40514 & w40504;
	assign w40511 = w40512 ^ w40514;
	assign w40501 = w40503 ^ w40511;
	assign w40505 = w40506 ^ w40514;
	assign w40491 = w40505 & w46252;
	assign w45071 = w40503 ^ w40521;
	assign w40495 = w45071 ^ w40473;
	assign w40484 = w40495 & w40536;
	assign w40493 = w40495 & w40532;
	assign w40462 = w46251 ^ w45071;
	assign w40502 = w40462 ^ w40425;
	assign w40492 = w40502 & w40531;
	assign w40483 = w40502 & w40533;
	assign w45070 = w40491 ^ w40493;
	assign w40510 = w40513 & w40511;
	assign w40421 = w40510 ^ w40522;
	assign w40417 = w40421 ^ w40457;
	assign w40416 = w46247 ^ w40417;
	assign w40420 = w46245 ^ w40417;
	assign w40497 = w40419 ^ w40420;
	assign w40509 = w40510 ^ w40472;
	assign w40500 = w40509 & w40501;
	assign w40423 = w40500 ^ w40524;
	assign w40415 = w40462 ^ w40423;
	assign w40494 = w40415 ^ w40416;
	assign w40465 = w40500 ^ w40475;
	assign w40499 = w40465 ^ w40467;
	assign w40422 = w40452 ^ w40415;
	assign w40498 = w40419 ^ w40422;
	assign w40418 = w40510 ^ w40466;
	assign w40496 = w40465 ^ w40418;
	assign w40486 = w40494 & w40527;
	assign w40480 = w40499 & w40534;
	assign w40487 = w40497 & w40529;
	assign w40443 = w40486 ^ w40487;
	assign w40489 = w40499 & w40538;
	assign w40447 = w40486 ^ w40489;
	assign w40444 = ~w40447;
	assign w40488 = w40509 & w40528;
	assign w40450 = w40488 ^ w40480;
	assign w40432 = w40488 ^ w40489;
	assign w40477 = w40494 & w40542;
	assign w40476 = w40498 & w40539;
	assign w40442 = w40487 ^ w40476;
	assign w40438 = ~w40442;
	assign w40485 = w40498 & w40530;
	assign w40479 = w40509 & w40535;
	assign w40481 = w40496 & w40541;
	assign w40463 = w40481 ^ w40485;
	assign w40441 = ~w40463;
	assign w40440 = w40441 ^ w40479;
	assign w40436 = w40440 ^ w45070;
	assign w50616 = w45213 ^ w9633;
	assign w46260 = w50616 ^ w480;
	assign w41128 = w46260 ^ w46254;
	assign w41198 = w41128 ^ w41123;
	assign w41208 = w46255 ^ w41128;
	assign w41204 = w46259 ^ w41208;
	assign w41207 = w46260 ^ w41083;
	assign w41193 = w46260 & w41207;
	assign w41191 = w41208 & w41204;
	assign w40482 = w40505 & w40537;
	assign w40478 = w40497 & w40540;
	assign w40439 = w40478 ^ w40436;
	assign w40543 = w40438 ^ w40439;
	assign w45068 = w40477 ^ w40478;
	assign w40459 = w40483 ^ w45068;
	assign w40460 = w40484 ^ w40459;
	assign w40435 = w40459 ^ w40436;
	assign w40464 = w40492 ^ w40460;
	assign w40469 = w40493 ^ w40464;
	assign w40433 = w40491 ^ w40464;
	assign w40544 = w40469 ^ w40443;
	assign w40446 = w40450 ^ w45068;
	assign w40449 = w45070 ^ w40446;
	assign w40445 = w40441 ^ w40446;
	assign w40545 = w40444 ^ w40445;
	assign w50875 = w40432 ^ w40433;
	assign w10198 = ~w50875;
	assign w50873 = ~w40545;
	assign w45838 = ~w40543;
	assign w45839 = ~w40544;
	assign w10321 = w45839 ^ w45838;
	assign w40490 = w40496 & w40526;
	assign w40448 = w40490 ^ w40481;
	assign w40546 = w40448 ^ w40449;
	assign w45069 = w40489 ^ w40490;
	assign w50876 = w45069 ^ w40469;
	assign w40471 = w40486 ^ w45069;
	assign w40437 = w40482 ^ w40471;
	assign w40434 = ~w40437;
	assign w50874 = w40434 ^ w40435;
	assign w40431 = w40487 ^ w40471;
	assign w50877 = w40460 ^ w40431;
	assign w45840 = ~w40546;
	assign w9579 = w50664 ^ w50654;
	assign w9915 = w9578 ^ w9579;
	assign w50524 = w9915 ^ w9880;
	assign w46352 = w50524 ^ w579;
	assign w41526 = w46352 ^ w46350;
	assign w41612 = w46352 ^ w46349;
	assign w41608 = w41612 ^ w41540;
	assign w41604 = w41523 ^ w41612;
	assign w41603 = w46356 ^ w41604;
	assign w41614 = w46354 ^ w46352;
	assign w41599 = w41524 ^ w41614;
	assign w41486 = w41526 ^ w41524;
	assign w41602 = w41523 ^ w41486;
	assign w41485 = w41526 ^ w46351;
	assign w41609 = w46356 ^ w41485;
	assign w41597 = w41604 & w41608;
	assign w41529 = w41597 ^ w41526;
	assign w41596 = w41605 & w41603;
	assign w41595 = w46356 & w41609;
	assign w41591 = w41612 & w41601;
	assign w41527 = w41591 ^ w41525;
	assign w41533 = w41529 ^ w41527;
	assign w41538 = w46349 ^ w41533;
	assign w41590 = w41614 & w41599;
	assign w41547 = w41590 ^ w41596;
	assign w41588 = w41547 ^ w41538;
	assign w41499 = w41590 ^ w41591;
	assign w41546 = w41499 ^ w41500;
	assign w41545 = w41546 ^ w41528;
	assign w41587 = w41593 ^ w41545;
	assign w41589 = w41611 & w41602;
	assign w41584 = w41588 & w41587;
	assign w45111 = w41589 ^ w41595;
	assign w41539 = w45111 ^ w41524;
	assign w41585 = w41547 ^ w41539;
	assign w41501 = w41533 ^ w45111;
	assign w41544 = w46351 ^ w41501;
	assign w41579 = w41584 ^ w41544;
	assign w45112 = w41589 ^ w41592;
	assign w41542 = w41590 ^ w45112;
	assign w41498 = w41593 ^ w41542;
	assign w41580 = w46355 ^ w41498;
	assign w41578 = w41579 & w41580;
	assign w41497 = w41578 ^ w41542;
	assign w41496 = w41578 ^ w41595;
	assign w41491 = w41496 ^ w41592;
	assign w41576 = w41584 ^ w41578;
	assign w41502 = w41528 ^ w45112;
	assign w41586 = w41502 ^ w41527;
	assign w41577 = w41578 ^ w41586;
	assign w41583 = w41584 ^ w41586;
	assign w41582 = w41585 & w41583;
	assign w41581 = w41582 ^ w41544;
	assign w41493 = w41582 ^ w41594;
	assign w41489 = w41493 ^ w41529;
	assign w41492 = w46349 ^ w41489;
	assign w41569 = w41491 ^ w41492;
	assign w41490 = w41582 ^ w41538;
	assign w41488 = w46351 ^ w41489;
	assign w41575 = w41586 & w41576;
	assign w41573 = w41575 ^ w41583;
	assign w41572 = w41581 & w41573;
	assign w41537 = w41572 ^ w41547;
	assign w41571 = w41537 ^ w41539;
	assign w41495 = w41572 ^ w41596;
	assign w41568 = w41537 ^ w41490;
	assign w41563 = w41577 & w46356;
	assign w41562 = w41568 & w41598;
	assign w41561 = w41571 & w41610;
	assign w41560 = w41581 & w41600;
	assign w41504 = w41560 ^ w41561;
	assign w41559 = w41569 & w41601;
	assign w41554 = w41577 & w41609;
	assign w41553 = w41568 & w41613;
	assign w41520 = w41562 ^ w41553;
	assign w41552 = w41571 & w41606;
	assign w41522 = w41560 ^ w41552;
	assign w41551 = w41581 & w41607;
	assign w41550 = w41569 & w41612;
	assign w45113 = w41561 ^ w41562;
	assign w45115 = w41575 ^ w41593;
	assign w41534 = w46355 ^ w45115;
	assign w41574 = w41534 ^ w41497;
	assign w41555 = w41574 & w41605;
	assign w41564 = w41574 & w41603;
	assign w41487 = w41534 ^ w41495;
	assign w41494 = w41524 ^ w41487;
	assign w41570 = w41491 ^ w41494;
	assign w41557 = w41570 & w41602;
	assign w41535 = w41553 ^ w41557;
	assign w41513 = ~w41535;
	assign w41512 = w41513 ^ w41551;
	assign w41566 = w41487 ^ w41488;
	assign w41549 = w41566 & w41614;
	assign w41548 = w41570 & w41611;
	assign w41514 = w41559 ^ w41548;
	assign w41510 = ~w41514;
	assign w43614 = w41549 ^ w41550;
	assign w41518 = w41522 ^ w43614;
	assign w41517 = w41513 ^ w41518;
	assign w41531 = w41555 ^ w43614;
	assign w41558 = w41566 & w41599;
	assign w41515 = w41558 ^ w41559;
	assign w41543 = w41558 ^ w45113;
	assign w41509 = w41554 ^ w41543;
	assign w41506 = ~w41509;
	assign w41503 = w41559 ^ w41543;
	assign w41519 = w41558 ^ w41561;
	assign w41516 = ~w41519;
	assign w41617 = w41516 ^ w41517;
	assign w41567 = w45115 ^ w41545;
	assign w41565 = w41567 & w41604;
	assign w41556 = w41567 & w41608;
	assign w41532 = w41556 ^ w41531;
	assign w41536 = w41564 ^ w41532;
	assign w41541 = w41565 ^ w41536;
	assign w50907 = w45113 ^ w41541;
	assign w41616 = w41541 ^ w41515;
	assign w41505 = w41563 ^ w41536;
	assign w50906 = w41504 ^ w41505;
	assign w50909 = w41532 ^ w41503;
	assign w50908 = ~w41616;
	assign w10241 = ~w50907;
	assign w45114 = w41563 ^ w41565;
	assign w41521 = w45114 ^ w41518;
	assign w41618 = w41520 ^ w41521;
	assign w41508 = w41512 ^ w45114;
	assign w41511 = w41550 ^ w41508;
	assign w41615 = w41510 ^ w41511;
	assign w41507 = w41531 ^ w41508;
	assign w50905 = w41506 ^ w41507;
	assign w45858 = ~w41617;
	assign w45859 = ~w41618;
	assign w45865 = ~w41615;
	assign w10414 = w41616 ^ w45865;
	assign w45950 = ~w9826;
	assign w9721 = w45950 ^ w50670;
	assign w50564 = w9720 ^ w9721;
	assign w9724 = w45950 ^ w50669;
	assign w50563 = w9723 ^ w9724;
	assign w46313 = w50563 ^ w554;
	assign w9728 = w45950 ^ w45872;
	assign w9726 = w9727 ^ w9728;
	assign w50561 = ~w9726;
	assign w46315 = w50561 ^ w552;
	assign w10174 = w46315 ^ w10178;
	assign w10161 = w10178 & w10174;
	assign w10091 = w46315 ^ w46313;
	assign w10108 = w46315 ^ w46314;
	assign w10173 = w10108 ^ w10175;
	assign w10068 = w46313 ^ w46314;
	assign w10181 = w46309 ^ w46315;
	assign w10093 = w46314 ^ w10091;
	assign w10168 = w10098 ^ w10093;
	assign w10160 = w10175 & w10168;
	assign w10169 = w46310 ^ w10093;
	assign w10166 = w46311 ^ w10093;
	assign w10162 = w10181 & w10166;
	assign w10096 = w10162 ^ w10092;
	assign w46312 = w50564 ^ w555;
	assign w10180 = w46312 ^ w46309;
	assign w10159 = w10180 & w10169;
	assign w10176 = w10180 ^ w10108;
	assign w10095 = w10159 ^ w10093;
	assign w10172 = w10091 ^ w10180;
	assign w10171 = w46316 ^ w10172;
	assign w10164 = w10173 & w10171;
	assign w10182 = w46314 ^ w46312;
	assign w10167 = w10092 ^ w10182;
	assign w10158 = w10182 & w10167;
	assign w10067 = w10158 ^ w10159;
	assign w10114 = w10067 ^ w10068;
	assign w10115 = w10158 ^ w10164;
	assign w10113 = w10114 ^ w10096;
	assign w10155 = w10161 ^ w10113;
	assign w10165 = w10172 & w10176;
	assign w10094 = w46312 ^ w46310;
	assign w10054 = w10094 ^ w10092;
	assign w10097 = w10165 ^ w10094;
	assign w10053 = w10094 ^ w46311;
	assign w10101 = w10097 ^ w10095;
	assign w10106 = w46309 ^ w10101;
	assign w10156 = w10115 ^ w10106;
	assign w10152 = w10156 & w10155;
	assign w10177 = w46316 ^ w10053;
	assign w10163 = w46316 & w10177;
	assign w10170 = w10091 ^ w10054;
	assign w10157 = w10179 & w10170;
	assign w43808 = w10157 ^ w10163;
	assign w10069 = w10101 ^ w43808;
	assign w10107 = w43808 ^ w10092;
	assign w10153 = w10115 ^ w10107;
	assign w10112 = w46311 ^ w10069;
	assign w10147 = w10152 ^ w10112;
	assign w43809 = w10157 ^ w10160;
	assign w10070 = w10096 ^ w43809;
	assign w10154 = w10070 ^ w10095;
	assign w10151 = w10152 ^ w10154;
	assign w10150 = w10153 & w10151;
	assign w10061 = w10150 ^ w10162;
	assign w10149 = w10150 ^ w10112;
	assign w10128 = w10149 & w10168;
	assign w10058 = w10150 ^ w10106;
	assign w10057 = w10061 ^ w10097;
	assign w10060 = w46309 ^ w10057;
	assign w10056 = w46311 ^ w10057;
	assign w10110 = w10158 ^ w43809;
	assign w10066 = w10161 ^ w10110;
	assign w10148 = w46315 ^ w10066;
	assign w10146 = w10147 & w10148;
	assign w10065 = w10146 ^ w10110;
	assign w10144 = w10152 ^ w10146;
	assign w10143 = w10154 & w10144;
	assign w43813 = w10143 ^ w10161;
	assign w10064 = w10146 ^ w10163;
	assign w10059 = w10064 ^ w10160;
	assign w10137 = w10059 ^ w10060;
	assign w10127 = w10137 & w10169;
	assign w10118 = w10137 & w10180;
	assign w10135 = w43813 ^ w10113;
	assign w10133 = w10135 & w10172;
	assign w10102 = w46315 ^ w43813;
	assign w10142 = w10102 ^ w10065;
	assign w10132 = w10142 & w10171;
	assign w10141 = w10143 ^ w10151;
	assign w10140 = w10149 & w10141;
	assign w10105 = w10140 ^ w10115;
	assign w10139 = w10105 ^ w10107;
	assign w10129 = w10139 & w10178;
	assign w10120 = w10139 & w10174;
	assign w10090 = w10128 ^ w10120;
	assign w10136 = w10105 ^ w10058;
	assign w10130 = w10136 & w10166;
	assign w43811 = w10129 ^ w10130;
	assign w10121 = w10136 & w10181;
	assign w10088 = w10130 ^ w10121;
	assign w10072 = w10128 ^ w10129;
	assign w10063 = w10140 ^ w10164;
	assign w10055 = w10102 ^ w10063;
	assign w10134 = w10055 ^ w10056;
	assign w10062 = w10092 ^ w10055;
	assign w10138 = w10059 ^ w10062;
	assign w10116 = w10138 & w10179;
	assign w10125 = w10138 & w10170;
	assign w10082 = w10127 ^ w10116;
	assign w10078 = ~w10082;
	assign w10117 = w10134 & w10182;
	assign w43810 = w10117 ^ w10118;
	assign w10086 = w10090 ^ w43810;
	assign w10103 = w10121 ^ w10125;
	assign w10081 = ~w10103;
	assign w10085 = w10081 ^ w10086;
	assign w10124 = w10135 & w10176;
	assign w10145 = w10146 ^ w10154;
	assign w10122 = w10145 & w10177;
	assign w10131 = w10145 & w46316;
	assign w43812 = w10131 ^ w10133;
	assign w10089 = w43812 ^ w10086;
	assign w10186 = w10088 ^ w10089;
	assign w45210 = ~w10186;
	assign w10498 = w45859 ^ w45210;
	assign w10123 = w10142 & w10173;
	assign w10099 = w10123 ^ w43810;
	assign w10100 = w10124 ^ w10099;
	assign w10104 = w10132 ^ w10100;
	assign w10109 = w10133 ^ w10104;
	assign w50912 = w43811 ^ w10109;
	assign w10501 = w50907 ^ w50912;
	assign w10073 = w10131 ^ w10104;
	assign w50911 = w10072 ^ w10073;
	assign w10240 = w50911 ^ w10241;
	assign w10119 = w10149 & w10175;
	assign w10080 = w10081 ^ w10119;
	assign w10076 = w10080 ^ w43812;
	assign w10079 = w10118 ^ w10076;
	assign w10075 = w10099 ^ w10076;
	assign w10183 = w10078 ^ w10079;
	assign w45212 = ~w10183;
	assign w10405 = w45212 ^ w50912;
	assign w10126 = w10134 & w10167;
	assign w10087 = w10126 ^ w10129;
	assign w10084 = ~w10087;
	assign w10185 = w10084 ^ w10085;
	assign w10111 = w10126 ^ w43811;
	assign w10077 = w10122 ^ w10111;
	assign w10074 = ~w10077;
	assign w50910 = w10074 ^ w10075;
	assign w10190 = w50911 ^ w50910;
	assign w10475 = w50905 ^ w50910;
	assign w10083 = w10126 ^ w10127;
	assign w10184 = w10109 ^ w10083;
	assign w45208 = ~w10184;
	assign w45209 = ~w10185;
	assign w10490 = w45858 ^ w45209;
	assign w10399 = ~w10490;
	assign w10071 = w10127 ^ w10111;
	assign w50913 = w10100 ^ w10071;
	assign w10436 = w50909 ^ w50913;
	assign w10427 = w50913 ^ w41616;
	assign w10500 = w50908 ^ w45208;
	assign w9754 = w45863 ^ w42822;
	assign w45952 = ~w9822;
	assign w9813 = w45952 ^ w45826;
	assign w50623 = w9813 ^ w9814;
	assign w9782 = w45952 ^ w50705;
	assign w9780 = w9781 ^ w9782;
	assign w9785 = w45952 ^ w45868;
	assign w50641 = w9784 ^ w9785;
	assign w50643 = ~w9780;
	assign w46233 = w50643 ^ w507;
	assign w38954 = w46233 ^ w46234;
	assign w46253 = w50623 ^ w487;
	assign w41211 = w46253 ^ w46259;
	assign w41209 = w46253 ^ w46258;
	assign w41192 = w41211 & w41196;
	assign w41122 = w46255 ^ w46253;
	assign w41084 = w41124 ^ w41122;
	assign w41205 = w41122 ^ w41128;
	assign w41190 = w41205 & w41198;
	assign w41200 = w41121 ^ w41084;
	assign w41187 = w41209 & w41200;
	assign w41197 = w41122 ^ w41212;
	assign w41188 = w41212 & w41197;
	assign w41210 = w46256 ^ w46253;
	assign w41202 = w41121 ^ w41210;
	assign w41189 = w41210 & w41199;
	assign w41097 = w41188 ^ w41189;
	assign w41144 = w41097 ^ w41098;
	assign w41206 = w41210 ^ w41138;
	assign w41195 = w41202 & w41206;
	assign w41127 = w41195 ^ w41124;
	assign w41201 = w46260 ^ w41202;
	assign w45094 = w41187 ^ w41193;
	assign w41137 = w45094 ^ w41122;
	assign w45095 = w41187 ^ w41190;
	assign w41140 = w41188 ^ w45095;
	assign w41096 = w41191 ^ w41140;
	assign w41178 = w46259 ^ w41096;
	assign w41203 = w41138 ^ w41205;
	assign w41194 = w41203 & w41201;
	assign w41125 = w41189 ^ w41123;
	assign w41131 = w41127 ^ w41125;
	assign w41136 = w46253 ^ w41131;
	assign w41099 = w41131 ^ w45094;
	assign w41142 = w46255 ^ w41099;
	assign w41145 = w41188 ^ w41194;
	assign w41186 = w41145 ^ w41136;
	assign w41183 = w41145 ^ w41137;
	assign w41126 = w41192 ^ w41122;
	assign w41143 = w41144 ^ w41126;
	assign w41100 = w41126 ^ w45095;
	assign w41184 = w41100 ^ w41125;
	assign w41185 = w41191 ^ w41143;
	assign w41182 = w41186 & w41185;
	assign w41181 = w41182 ^ w41184;
	assign w41180 = w41183 & w41181;
	assign w41088 = w41180 ^ w41136;
	assign w41091 = w41180 ^ w41192;
	assign w41087 = w41091 ^ w41127;
	assign w41090 = w46253 ^ w41087;
	assign w41086 = w46255 ^ w41087;
	assign w41177 = w41182 ^ w41142;
	assign w41176 = w41177 & w41178;
	assign w41094 = w41176 ^ w41193;
	assign w41095 = w41176 ^ w41140;
	assign w41089 = w41094 ^ w41190;
	assign w41167 = w41089 ^ w41090;
	assign w41148 = w41167 & w41210;
	assign w41157 = w41167 & w41199;
	assign w41175 = w41176 ^ w41184;
	assign w41161 = w41175 & w46260;
	assign w41152 = w41175 & w41207;
	assign w41174 = w41182 ^ w41176;
	assign w41173 = w41184 & w41174;
	assign w41171 = w41173 ^ w41181;
	assign w41179 = w41180 ^ w41142;
	assign w41158 = w41179 & w41198;
	assign w41149 = w41179 & w41205;
	assign w41170 = w41179 & w41171;
	assign w41135 = w41170 ^ w41145;
	assign w41166 = w41135 ^ w41088;
	assign w41151 = w41166 & w41211;
	assign w41160 = w41166 & w41196;
	assign w41093 = w41170 ^ w41194;
	assign w41118 = w41160 ^ w41151;
	assign w41169 = w41135 ^ w41137;
	assign w41159 = w41169 & w41208;
	assign w41150 = w41169 & w41204;
	assign w41120 = w41158 ^ w41150;
	assign w41102 = w41158 ^ w41159;
	assign w45097 = w41159 ^ w41160;
	assign w45099 = w41173 ^ w41191;
	assign w41132 = w46259 ^ w45099;
	assign w41172 = w41132 ^ w41095;
	assign w41162 = w41172 & w41201;
	assign w41153 = w41172 & w41203;
	assign w41085 = w41132 ^ w41093;
	assign w41092 = w41122 ^ w41085;
	assign w41168 = w41089 ^ w41092;
	assign w41146 = w41168 & w41209;
	assign w41112 = w41157 ^ w41146;
	assign w41164 = w41085 ^ w41086;
	assign w41156 = w41164 & w41197;
	assign w41113 = w41156 ^ w41157;
	assign w41117 = w41156 ^ w41159;
	assign w41114 = ~w41117;
	assign w41155 = w41168 & w41200;
	assign w41141 = w41156 ^ w45097;
	assign w41147 = w41164 & w41212;
	assign w41107 = w41152 ^ w41141;
	assign w41104 = ~w41107;
	assign w41133 = w41151 ^ w41155;
	assign w41111 = ~w41133;
	assign w41110 = w41111 ^ w41149;
	assign w41108 = ~w41112;
	assign w41101 = w41157 ^ w41141;
	assign w41165 = w45099 ^ w41143;
	assign w41154 = w41165 & w41206;
	assign w41163 = w41165 & w41202;
	assign w45096 = w41147 ^ w41148;
	assign w41116 = w41120 ^ w45096;
	assign w41115 = w41111 ^ w41116;
	assign w41215 = w41114 ^ w41115;
	assign w41129 = w41153 ^ w45096;
	assign w41130 = w41154 ^ w41129;
	assign w50889 = w41130 ^ w41101;
	assign w41134 = w41162 ^ w41130;
	assign w41139 = w41163 ^ w41134;
	assign w41214 = w41139 ^ w41113;
	assign w50888 = w45097 ^ w41139;
	assign w41103 = w41161 ^ w41134;
	assign w50887 = w41102 ^ w41103;
	assign w45846 = ~w41215;
	assign w45853 = ~w41214;
	assign w46235 = w50641 ^ w505;
	assign w38977 = w46235 ^ w46233;
	assign w38979 = w46234 ^ w38977;
	assign w39052 = w46231 ^ w38979;
	assign w39054 = w38984 ^ w38979;
	assign w39060 = w46235 ^ w39064;
	assign w39055 = w46230 ^ w38979;
	assign w39056 = w38977 ^ w38940;
	assign w39043 = w39065 & w39056;
	assign w39046 = w39061 & w39054;
	assign w39047 = w39064 & w39060;
	assign w39058 = w38977 ^ w39066;
	assign w39057 = w46236 ^ w39058;
	assign w38994 = w46235 ^ w46234;
	assign w39059 = w38994 ^ w39061;
	assign w39050 = w39059 & w39057;
	assign w39062 = w39066 ^ w38994;
	assign w39001 = w39044 ^ w39050;
	assign w39045 = w39066 & w39055;
	assign w38981 = w39045 ^ w38979;
	assign w38953 = w39044 ^ w39045;
	assign w39067 = w46229 ^ w46235;
	assign w39048 = w39067 & w39052;
	assign w38982 = w39048 ^ w38978;
	assign w39051 = w39058 & w39062;
	assign w38983 = w39051 ^ w38980;
	assign w45004 = w39043 ^ w39046;
	assign w38956 = w38982 ^ w45004;
	assign w39040 = w38956 ^ w38981;
	assign w38996 = w39044 ^ w45004;
	assign w45007 = w39043 ^ w39049;
	assign w38993 = w45007 ^ w38978;
	assign w39039 = w39001 ^ w38993;
	assign w38987 = w38983 ^ w38981;
	assign w38955 = w38987 ^ w45007;
	assign w38998 = w46231 ^ w38955;
	assign w38992 = w46229 ^ w38987;
	assign w39042 = w39001 ^ w38992;
	assign w39000 = w38953 ^ w38954;
	assign w38999 = w39000 ^ w38982;
	assign w39041 = w39047 ^ w38999;
	assign w39038 = w39042 & w39041;
	assign w39033 = w39038 ^ w38998;
	assign w39037 = w39038 ^ w39040;
	assign w39036 = w39039 & w39037;
	assign w39035 = w39036 ^ w38998;
	assign w38944 = w39036 ^ w38992;
	assign w39014 = w39035 & w39054;
	assign w39005 = w39035 & w39061;
	assign w38947 = w39036 ^ w39048;
	assign w38943 = w38947 ^ w38983;
	assign w38942 = w46231 ^ w38943;
	assign w38946 = w46229 ^ w38943;
	assign w38952 = w39047 ^ w38996;
	assign w39034 = w46235 ^ w38952;
	assign w39032 = w39033 & w39034;
	assign w39031 = w39032 ^ w39040;
	assign w39030 = w39038 ^ w39032;
	assign w38951 = w39032 ^ w38996;
	assign w38950 = w39032 ^ w39049;
	assign w39029 = w39040 & w39030;
	assign w39027 = w39029 ^ w39037;
	assign w39026 = w39035 & w39027;
	assign w39008 = w39031 & w39063;
	assign w38949 = w39026 ^ w39050;
	assign w38991 = w39026 ^ w39001;
	assign w39025 = w38991 ^ w38993;
	assign w39015 = w39025 & w39064;
	assign w38958 = w39014 ^ w39015;
	assign w39017 = w39031 & w46236;
	assign w45006 = w39029 ^ w39047;
	assign w39021 = w45006 ^ w38999;
	assign w39010 = w39021 & w39062;
	assign w39019 = w39021 & w39058;
	assign w45009 = w39017 ^ w39019;
	assign w38988 = w46235 ^ w45006;
	assign w38941 = w38988 ^ w38949;
	assign w39028 = w38988 ^ w38951;
	assign w39020 = w38941 ^ w38942;
	assign w39009 = w39028 & w39059;
	assign w39018 = w39028 & w39057;
	assign w39012 = w39020 & w39053;
	assign w38973 = w39012 ^ w39015;
	assign w38970 = ~w38973;
	assign w38948 = w38978 ^ w38941;
	assign w39022 = w38991 ^ w38944;
	assign w39007 = w39022 & w39067;
	assign w39016 = w39022 & w39052;
	assign w38974 = w39016 ^ w39007;
	assign w45008 = w39015 ^ w39016;
	assign w38997 = w39012 ^ w45008;
	assign w38963 = w39008 ^ w38997;
	assign w38960 = ~w38963;
	assign w38945 = w38950 ^ w39046;
	assign w39023 = w38945 ^ w38946;
	assign w39004 = w39023 & w39066;
	assign w39024 = w38945 ^ w38948;
	assign w39002 = w39024 & w39065;
	assign w39011 = w39024 & w39056;
	assign w38989 = w39007 ^ w39011;
	assign w38967 = ~w38989;
	assign w38966 = w38967 ^ w39005;
	assign w38962 = w38966 ^ w45009;
	assign w39013 = w39023 & w39055;
	assign w38969 = w39012 ^ w39013;
	assign w38957 = w39013 ^ w38997;
	assign w38968 = w39013 ^ w39002;
	assign w38964 = ~w38968;
	assign w38965 = w39004 ^ w38962;
	assign w39069 = w38964 ^ w38965;
	assign w39006 = w39025 & w39060;
	assign w38976 = w39014 ^ w39006;
	assign w39003 = w39020 & w39068;
	assign w45005 = w39003 ^ w39004;
	assign w38972 = w38976 ^ w45005;
	assign w38975 = w45009 ^ w38972;
	assign w39072 = w38974 ^ w38975;
	assign w38971 = w38967 ^ w38972;
	assign w39071 = w38970 ^ w38971;
	assign w38985 = w39009 ^ w45005;
	assign w38986 = w39010 ^ w38985;
	assign w38990 = w39018 ^ w38986;
	assign w38959 = w39017 ^ w38990;
	assign w38995 = w39019 ^ w38990;
	assign w39070 = w38995 ^ w38969;
	assign w50921 = w38986 ^ w38957;
	assign w50919 = w38958 ^ w38959;
	assign w10461 = w50906 ^ w50919;
	assign w10420 = w10475 ^ w10461;
	assign w10418 = ~w10420;
	assign w38961 = w38985 ^ w38962;
	assign w50920 = w45008 ^ w38995;
	assign w10430 = w50920 ^ w10241;
	assign w10401 = w10436 ^ w50921;
	assign w50918 = w38960 ^ w38961;
	assign w10408 = w10475 ^ w50918;
	assign w10204 = w50919 ^ w50918;
	assign w10447 = w50909 ^ w50921;
	assign w10203 = w10447 ^ w50905;
	assign w10523 = w10203 ^ w10204;
	assign w10201 = w10447 ^ w45859;
	assign w10433 = w10447 ^ w50912;
	assign w45802 = ~w39071;
	assign w10245 = w45802 ^ w50910;
	assign w45803 = ~w39072;
	assign w10202 = w45803 ^ w45209;
	assign w10524 = w10201 ^ w10202;
	assign w45808 = ~w39069;
	assign w10390 = w10500 ^ w45808;
	assign w10470 = w45865 ^ w45808;
	assign w10417 = w10501 ^ w10470;
	assign w45809 = ~w39070;
	assign w45098 = w41161 ^ w41163;
	assign w41106 = w41110 ^ w45098;
	assign w41109 = w41148 ^ w41106;
	assign w41105 = w41129 ^ w41106;
	assign w50886 = w41104 ^ w41105;
	assign w41213 = w41108 ^ w41109;
	assign w45852 = ~w41213;
	assign w41119 = w45098 ^ w41116;
	assign w41216 = w41118 ^ w41119;
	assign w45847 = ~w41216;
	assign w45953 = ~w9829;
	assign w9753 = w45953 ^ w50667;
	assign w50543 = w9753 ^ w9754;
	assign w46333 = w50543 ^ w598;
	assign w42596 = w46335 ^ w46333;
	assign w42679 = w42596 ^ w42602;
	assign w42677 = w42612 ^ w42679;
	assign w42685 = w46333 ^ w46339;
	assign w42683 = w46333 ^ w46338;
	assign w42666 = w42685 & w42670;
	assign w42600 = w42666 ^ w42596;
	assign w42664 = w42679 & w42672;
	assign w9617 = w45953 ^ w45882;
	assign w9899 = w9617 ^ w9618;
	assign w50529 = w9899 ^ w9891;
	assign w46347 = w50529 ^ w584;
	assign w40809 = w46341 ^ w46347;
	assign w40736 = w46347 ^ w46346;
	assign w40801 = w40736 ^ w40803;
	assign w40802 = w46347 ^ w40806;
	assign w40719 = w46347 ^ w46345;
	assign w9774 = w45953 ^ w50650;
	assign w50532 = w9773 ^ w9774;
	assign w46344 = w50532 ^ w587;
	assign w40808 = w46344 ^ w46341;
	assign w40804 = w40808 ^ w40736;
	assign w40800 = w40719 ^ w40808;
	assign w40722 = w46344 ^ w46342;
	assign w40682 = w40722 ^ w40720;
	assign w40798 = w40719 ^ w40682;
	assign w40681 = w40722 ^ w46343;
	assign w40805 = w46348 ^ w40681;
	assign w40799 = w46348 ^ w40800;
	assign w40793 = w40800 & w40804;
	assign w40725 = w40793 ^ w40722;
	assign w40792 = w40801 & w40799;
	assign w40785 = w40807 & w40798;
	assign w40810 = w46346 ^ w46344;
	assign w40795 = w40720 ^ w40810;
	assign w40786 = w40810 & w40795;
	assign w40791 = w46348 & w40805;
	assign w40743 = w40786 ^ w40792;
	assign w40721 = w46346 ^ w40719;
	assign w40797 = w46342 ^ w40721;
	assign w40794 = w46343 ^ w40721;
	assign w40796 = w40726 ^ w40721;
	assign w40788 = w40803 & w40796;
	assign w40790 = w40809 & w40794;
	assign w40724 = w40790 ^ w40720;
	assign w40787 = w40808 & w40797;
	assign w40723 = w40787 ^ w40721;
	assign w40729 = w40725 ^ w40723;
	assign w40734 = w46341 ^ w40729;
	assign w40784 = w40743 ^ w40734;
	assign w45078 = w40785 ^ w40788;
	assign w40698 = w40724 ^ w45078;
	assign w40782 = w40698 ^ w40723;
	assign w40738 = w40786 ^ w45078;
	assign w40695 = w40786 ^ w40787;
	assign w40742 = w40695 ^ w40696;
	assign w40741 = w40742 ^ w40724;
	assign w40789 = w40806 & w40802;
	assign w40783 = w40789 ^ w40741;
	assign w40694 = w40789 ^ w40738;
	assign w40776 = w46347 ^ w40694;
	assign w40780 = w40784 & w40783;
	assign w40779 = w40780 ^ w40782;
	assign w45077 = w40785 ^ w40791;
	assign w40735 = w45077 ^ w40720;
	assign w40781 = w40743 ^ w40735;
	assign w40778 = w40781 & w40779;
	assign w40689 = w40778 ^ w40790;
	assign w40685 = w40689 ^ w40725;
	assign w40688 = w46341 ^ w40685;
	assign w40684 = w46343 ^ w40685;
	assign w40686 = w40778 ^ w40734;
	assign w40697 = w40729 ^ w45077;
	assign w40740 = w46343 ^ w40697;
	assign w40775 = w40780 ^ w40740;
	assign w40774 = w40775 & w40776;
	assign w40772 = w40780 ^ w40774;
	assign w40771 = w40782 & w40772;
	assign w40692 = w40774 ^ w40791;
	assign w40687 = w40692 ^ w40788;
	assign w40765 = w40687 ^ w40688;
	assign w40746 = w40765 & w40808;
	assign w40769 = w40771 ^ w40779;
	assign w40693 = w40774 ^ w40738;
	assign w40755 = w40765 & w40797;
	assign w40773 = w40774 ^ w40782;
	assign w40750 = w40773 & w40805;
	assign w40759 = w40773 & w46348;
	assign w45082 = w40771 ^ w40789;
	assign w40730 = w46347 ^ w45082;
	assign w40770 = w40730 ^ w40693;
	assign w40760 = w40770 & w40799;
	assign w40751 = w40770 & w40801;
	assign w40763 = w45082 ^ w40741;
	assign w40761 = w40763 & w40800;
	assign w40752 = w40763 & w40804;
	assign w40777 = w40778 ^ w40740;
	assign w40768 = w40777 & w40769;
	assign w40733 = w40768 ^ w40743;
	assign w40764 = w40733 ^ w40686;
	assign w40756 = w40777 & w40796;
	assign w40767 = w40733 ^ w40735;
	assign w40757 = w40767 & w40806;
	assign w40700 = w40756 ^ w40757;
	assign w40749 = w40764 & w40809;
	assign w40691 = w40768 ^ w40792;
	assign w40683 = w40730 ^ w40691;
	assign w40690 = w40720 ^ w40683;
	assign w40766 = w40687 ^ w40690;
	assign w40744 = w40766 & w40807;
	assign w40762 = w40683 ^ w40684;
	assign w40754 = w40762 & w40795;
	assign w40715 = w40754 ^ w40757;
	assign w40712 = ~w40715;
	assign w40711 = w40754 ^ w40755;
	assign w40747 = w40777 & w40803;
	assign w40753 = w40766 & w40798;
	assign w40731 = w40749 ^ w40753;
	assign w40709 = ~w40731;
	assign w40708 = w40709 ^ w40747;
	assign w40745 = w40762 & w40810;
	assign w45079 = w40745 ^ w40746;
	assign w40727 = w40751 ^ w45079;
	assign w40728 = w40752 ^ w40727;
	assign w40732 = w40760 ^ w40728;
	assign w40701 = w40759 ^ w40732;
	assign w50892 = w40700 ^ w40701;
	assign w10217 = ~w50892;
	assign w10227 = w50898 ^ w10217;
	assign w10216 = w10217 ^ w50886;
	assign w40758 = w40764 & w40794;
	assign w45080 = w40757 ^ w40758;
	assign w10488 = w50887 ^ w50892;
	assign w10255 = ~w10488;
	assign w40748 = w40767 & w40802;
	assign w40718 = w40756 ^ w40748;
	assign w40714 = w40718 ^ w45079;
	assign w40713 = w40709 ^ w40714;
	assign w40813 = w40712 ^ w40713;
	assign w50890 = ~w40813;
	assign w10502 = w45846 ^ w50890;
	assign w10270 = w45854 ^ w40813;
	assign w10213 = w40813 ^ w45847;
	assign w40710 = w40755 ^ w40744;
	assign w40706 = ~w40710;
	assign w40716 = w40758 ^ w40749;
	assign w40739 = w40754 ^ w45080;
	assign w40705 = w40750 ^ w40739;
	assign w40702 = ~w40705;
	assign w40699 = w40755 ^ w40739;
	assign w50896 = w40728 ^ w40699;
	assign w10288 = w50896 ^ w45853;
	assign w10444 = w50896 ^ w50900;
	assign w10225 = ~w10444;
	assign w10440 = w50889 ^ w50896;
	assign w45894 = ~w10440;
	assign w10279 = w45894 ^ w50888;
	assign w10281 = w45894 ^ w50887;
	assign w10285 = w45894 ^ w45846;
	assign w45081 = w40759 ^ w40761;
	assign w40704 = w40708 ^ w45081;
	assign w40703 = w40727 ^ w40704;
	assign w40707 = w40746 ^ w40704;
	assign w40811 = w40706 ^ w40707;
	assign w10265 = w45860 ^ w40811;
	assign w50894 = ~w40811;
	assign w10473 = w45852 ^ w50894;
	assign w10296 = w40811 ^ w50888;
	assign w50891 = w40702 ^ w40703;
	assign w10224 = ~w50891;
	assign w10299 = w10224 ^ w45846;
	assign w10223 = w50897 ^ w10224;
	assign w10495 = w50886 ^ w50891;
	assign w10271 = ~w10495;
	assign w40717 = w45081 ^ w40714;
	assign w40814 = w40716 ^ w40717;
	assign w45843 = ~w40814;
	assign w10503 = w45847 ^ w45843;
	assign w10272 = w10503 ^ w10444;
	assign w10221 = w45855 ^ w45843;
	assign w40737 = w40761 ^ w40732;
	assign w50893 = w45080 ^ w40737;
	assign w10480 = w50888 ^ w50893;
	assign w10268 = w50899 ^ w50893;
	assign w40812 = w40737 ^ w40711;
	assign w50895 = ~w40812;
	assign w10466 = w45853 ^ w50895;
	assign w10263 = w45861 ^ w40812;
	assign w10291 = w40812 ^ w45852;
	assign w10252 = ~w10480;
	assign w10219 = w50893 ^ w50887;
	assign w45959 = ~w10436;
	assign w10239 = w45959 ^ w50906;
	assign w10508 = w10239 ^ w10240;
	assign w10424 = w45959 ^ w45858;
	assign w45961 = ~w43075;
	assign w42897 = w45961 ^ w45301;
	assign w50408 = w42896 ^ w42897;
	assign w42892 = w45961 ^ w50496;
	assign w50410 = w42891 ^ w42892;
	assign w42889 = w45961 ^ w50497;
	assign w50411 = w42888 ^ w42889;
	assign w46393 = w50410 ^ w411;
	assign w46395 = w50408 ^ w409;
	assign w39396 = w46395 ^ w46394;
	assign w39461 = w39396 ^ w39463;
	assign w46392 = w50411 ^ w412;
	assign w39468 = w46392 ^ w46389;
	assign w39464 = w39468 ^ w39396;
	assign w39470 = w46394 ^ w46392;
	assign w39455 = w39380 ^ w39470;
	assign w39462 = w46395 ^ w39466;
	assign w39449 = w39466 & w39462;
	assign w39379 = w46395 ^ w46393;
	assign w39381 = w46394 ^ w39379;
	assign w39457 = w46390 ^ w39381;
	assign w39460 = w39379 ^ w39468;
	assign w39459 = w46396 ^ w39460;
	assign w39456 = w39386 ^ w39381;
	assign w39447 = w39468 & w39457;
	assign w39383 = w39447 ^ w39381;
	assign w39448 = w39463 & w39456;
	assign w39356 = w46393 ^ w46394;
	assign w39446 = w39470 & w39455;
	assign w39355 = w39446 ^ w39447;
	assign w39402 = w39355 ^ w39356;
	assign w39453 = w39460 & w39464;
	assign w39382 = w46392 ^ w46390;
	assign w39342 = w39382 ^ w39380;
	assign w39385 = w39453 ^ w39382;
	assign w39389 = w39385 ^ w39383;
	assign w39394 = w46389 ^ w39389;
	assign w39458 = w39379 ^ w39342;
	assign w39341 = w39382 ^ w46391;
	assign w39465 = w46396 ^ w39341;
	assign w39469 = w46389 ^ w46395;
	assign w39452 = w39461 & w39459;
	assign w39403 = w39446 ^ w39452;
	assign w39444 = w39403 ^ w39394;
	assign w39451 = w46396 & w39465;
	assign w39454 = w46391 ^ w39381;
	assign w39450 = w39469 & w39454;
	assign w39384 = w39450 ^ w39380;
	assign w39401 = w39402 ^ w39384;
	assign w39443 = w39449 ^ w39401;
	assign w39440 = w39444 & w39443;
	assign w39221 = w39312 ^ w39313;
	assign w39268 = w39221 ^ w39222;
	assign w39267 = w39268 ^ w39250;
	assign w39309 = w39315 ^ w39267;
	assign w39306 = w39310 & w39309;
	assign w39301 = w39306 ^ w39266;
	assign w39300 = w39301 & w39302;
	assign w39219 = w39300 ^ w39264;
	assign w39299 = w39300 ^ w39308;
	assign w39218 = w39300 ^ w39317;
	assign w39285 = w39299 & w46332;
	assign w39213 = w39218 ^ w39314;
	assign w39276 = w39299 & w39331;
	assign w39305 = w39306 ^ w39308;
	assign w39304 = w39307 & w39305;
	assign w39303 = w39304 ^ w39266;
	assign w39282 = w39303 & w39322;
	assign w39215 = w39304 ^ w39316;
	assign w39211 = w39215 ^ w39251;
	assign w39273 = w39303 & w39329;
	assign w39212 = w39304 ^ w39260;
	assign w39214 = w46325 ^ w39211;
	assign w39291 = w39213 ^ w39214;
	assign w39272 = w39291 & w39334;
	assign w39281 = w39291 & w39323;
	assign w39210 = w46327 ^ w39211;
	assign w39298 = w39306 ^ w39300;
	assign w39297 = w39308 & w39298;
	assign w45020 = w39297 ^ w39315;
	assign w39289 = w45020 ^ w39267;
	assign w39287 = w39289 & w39326;
	assign w39278 = w39289 & w39330;
	assign w45019 = w39285 ^ w39287;
	assign w39256 = w46331 ^ w45020;
	assign w39296 = w39256 ^ w39219;
	assign w39277 = w39296 & w39327;
	assign w39286 = w39296 & w39325;
	assign w39295 = w39297 ^ w39305;
	assign w39294 = w39303 & w39295;
	assign w39217 = w39294 ^ w39318;
	assign w39209 = w39256 ^ w39217;
	assign w39216 = w39246 ^ w39209;
	assign w39292 = w39213 ^ w39216;
	assign w39270 = w39292 & w39333;
	assign w39236 = w39281 ^ w39270;
	assign w39288 = w39209 ^ w39210;
	assign w39271 = w39288 & w39336;
	assign w39279 = w39292 & w39324;
	assign w39232 = ~w39236;
	assign w45017 = w39271 ^ w39272;
	assign w39253 = w39277 ^ w45017;
	assign w39280 = w39288 & w39321;
	assign w39237 = w39280 ^ w39281;
	assign w39254 = w39278 ^ w39253;
	assign w39258 = w39286 ^ w39254;
	assign w39227 = w39285 ^ w39258;
	assign w39263 = w39287 ^ w39258;
	assign w39259 = w39294 ^ w39269;
	assign w39293 = w39259 ^ w39261;
	assign w39290 = w39259 ^ w39212;
	assign w39274 = w39293 & w39328;
	assign w39244 = w39282 ^ w39274;
	assign w39240 = w39244 ^ w45017;
	assign w39243 = w45019 ^ w39240;
	assign w39275 = w39290 & w39335;
	assign w39284 = w39290 & w39320;
	assign w39283 = w39293 & w39332;
	assign w39226 = w39282 ^ w39283;
	assign w39241 = w39280 ^ w39283;
	assign w39238 = ~w39241;
	assign w50865 = w39226 ^ w39227;
	assign w39257 = w39275 ^ w39279;
	assign w39235 = ~w39257;
	assign w39234 = w39235 ^ w39273;
	assign w45018 = w39283 ^ w39284;
	assign w50866 = w45018 ^ w39263;
	assign w10493 = w50862 ^ w50866;
	assign w39265 = w39280 ^ w45018;
	assign w10496 = w50861 ^ w50865;
	assign w39242 = w39284 ^ w39275;
	assign w39340 = w39242 ^ w39243;
	assign w45811 = ~w39340;
	assign w39239 = w39235 ^ w39240;
	assign w39339 = w39238 ^ w39239;
	assign w45810 = ~w39339;
	assign w10363 = w45810 ^ w42421;
	assign w39338 = w39263 ^ w39237;
	assign w50867 = ~w39338;
	assign w10486 = w45876 ^ w50867;
	assign w39230 = w39234 ^ w45019;
	assign w39233 = w39272 ^ w39230;
	assign w39337 = w39232 ^ w39233;
	assign w39229 = w39253 ^ w39230;
	assign w45817 = ~w39337;
	assign w10489 = w45875 ^ w45817;
	assign w39231 = w39276 ^ w39265;
	assign w39228 = ~w39231;
	assign w50864 = w39228 ^ w39229;
	assign w39225 = w39281 ^ w39265;
	assign w50868 = w39254 ^ w39225;
	assign w10441 = w50863 ^ w50868;
	assign w10234 = w10441 ^ w45811;
	assign w45956 = ~w10441;
	assign w10236 = w45956 ^ w50864;
	assign w10509 = w10236 ^ w10237;
	assign w10360 = w45956 ^ w50862;
	assign w39445 = w39467 & w39458;
	assign w45021 = w39445 ^ w39448;
	assign w45024 = w39445 ^ w39451;
	assign w39395 = w45024 ^ w39380;
	assign w39441 = w39403 ^ w39395;
	assign w39398 = w39446 ^ w45021;
	assign w39357 = w39389 ^ w45024;
	assign w39400 = w46391 ^ w39357;
	assign w39435 = w39440 ^ w39400;
	assign w39358 = w39384 ^ w45021;
	assign w39442 = w39358 ^ w39383;
	assign w39439 = w39440 ^ w39442;
	assign w39354 = w39449 ^ w39398;
	assign w39436 = w46395 ^ w39354;
	assign w39434 = w39435 & w39436;
	assign w39352 = w39434 ^ w39451;
	assign w39347 = w39352 ^ w39448;
	assign w39353 = w39434 ^ w39398;
	assign w39433 = w39434 ^ w39442;
	assign w39419 = w39433 & w46396;
	assign w39410 = w39433 & w39465;
	assign w39432 = w39440 ^ w39434;
	assign w39431 = w39442 & w39432;
	assign w45023 = w39431 ^ w39449;
	assign w39390 = w46395 ^ w45023;
	assign w39430 = w39390 ^ w39353;
	assign w39420 = w39430 & w39459;
	assign w39411 = w39430 & w39461;
	assign w39429 = w39431 ^ w39439;
	assign w39423 = w45023 ^ w39401;
	assign w39421 = w39423 & w39460;
	assign w39412 = w39423 & w39464;
	assign w45026 = w39419 ^ w39421;
	assign w46322 = w50554 ^ w545;
	assign w9959 = w46322 ^ w9957;
	assign w10032 = w46319 ^ w9959;
	assign w10035 = w46318 ^ w9959;
	assign w10048 = w46322 ^ w46320;
	assign w10033 = w9958 ^ w10048;
	assign w10034 = w9964 ^ w9959;
	assign w9934 = w46321 ^ w46322;
	assign w10025 = w10046 & w10035;
	assign w9961 = w10025 ^ w9959;
	assign w10026 = w10041 & w10034;
	assign w10045 = w46317 ^ w46322;
	assign w10023 = w10045 & w10036;
	assign w43804 = w10023 ^ w10026;
	assign w43803 = w10023 ^ w10029;
	assign w9973 = w43803 ^ w9958;
	assign w9974 = w46323 ^ w46322;
	assign w10039 = w9974 ^ w10041;
	assign w10030 = w10039 & w10037;
	assign w10042 = w10046 ^ w9974;
	assign w10031 = w10038 & w10042;
	assign w9963 = w10031 ^ w9960;
	assign w9967 = w9963 ^ w9961;
	assign w9972 = w46317 ^ w9967;
	assign w9935 = w9967 ^ w43803;
	assign w9978 = w46319 ^ w9935;
	assign w10024 = w10048 & w10033;
	assign w9933 = w10024 ^ w10025;
	assign w9980 = w9933 ^ w9934;
	assign w9976 = w10024 ^ w43804;
	assign w9932 = w10027 ^ w9976;
	assign w10014 = w46323 ^ w9932;
	assign w9981 = w10024 ^ w10030;
	assign w10019 = w9981 ^ w9973;
	assign w10022 = w9981 ^ w9972;
	assign w10028 = w10047 & w10032;
	assign w9962 = w10028 ^ w9958;
	assign w9979 = w9980 ^ w9962;
	assign w9936 = w9962 ^ w43804;
	assign w10020 = w9936 ^ w9961;
	assign w10021 = w10027 ^ w9979;
	assign w10018 = w10022 & w10021;
	assign w10017 = w10018 ^ w10020;
	assign w10016 = w10019 & w10017;
	assign w10013 = w10018 ^ w9978;
	assign w10012 = w10013 & w10014;
	assign w10011 = w10012 ^ w10020;
	assign w9930 = w10012 ^ w10029;
	assign w9925 = w9930 ^ w10026;
	assign w9931 = w10012 ^ w9976;
	assign w9927 = w10016 ^ w10028;
	assign w9923 = w9927 ^ w9963;
	assign w9926 = w46317 ^ w9923;
	assign w10003 = w9925 ^ w9926;
	assign w9984 = w10003 & w10046;
	assign w9924 = w10016 ^ w9972;
	assign w10010 = w10018 ^ w10012;
	assign w10009 = w10020 & w10010;
	assign w10007 = w10009 ^ w10017;
	assign w10015 = w10016 ^ w9978;
	assign w9994 = w10015 & w10034;
	assign w9985 = w10015 & w10041;
	assign w10006 = w10015 & w10007;
	assign w9929 = w10006 ^ w10030;
	assign w9971 = w10006 ^ w9981;
	assign w10005 = w9971 ^ w9973;
	assign w9986 = w10005 & w10040;
	assign w9956 = w9994 ^ w9986;
	assign w9995 = w10005 & w10044;
	assign w9938 = w9994 ^ w9995;
	assign w10002 = w9971 ^ w9924;
	assign w9996 = w10002 & w10032;
	assign w43805 = w9995 ^ w9996;
	assign w9987 = w10002 & w10047;
	assign w9954 = w9996 ^ w9987;
	assign w9993 = w10003 & w10035;
	assign w9988 = w10011 & w10043;
	assign w9922 = w46319 ^ w9923;
	assign w43807 = w10009 ^ w10027;
	assign w10001 = w43807 ^ w9979;
	assign w9999 = w10001 & w10038;
	assign w9990 = w10001 & w10042;
	assign w9968 = w46323 ^ w43807;
	assign w9921 = w9968 ^ w9929;
	assign w10000 = w9921 ^ w9922;
	assign w9983 = w10000 & w10048;
	assign w43524 = w9983 ^ w9984;
	assign w9952 = w9956 ^ w43524;
	assign w9992 = w10000 & w10033;
	assign w9953 = w9992 ^ w9995;
	assign w9949 = w9992 ^ w9993;
	assign w10008 = w9968 ^ w9931;
	assign w9989 = w10008 & w10039;
	assign w9965 = w9989 ^ w43524;
	assign w9966 = w9990 ^ w9965;
	assign w9998 = w10008 & w10037;
	assign w9950 = ~w9953;
	assign w9970 = w9998 ^ w9966;
	assign w9975 = w9999 ^ w9970;
	assign w10050 = w9975 ^ w9949;
	assign w50851 = w43805 ^ w9975;
	assign w45205 = ~w10050;
	assign w9977 = w9992 ^ w43805;
	assign w9937 = w9993 ^ w9977;
	assign w9943 = w9988 ^ w9977;
	assign w9940 = ~w9943;
	assign w50852 = w9966 ^ w9937;
	assign w10312 = w10489 ^ w50851;
	assign w10310 = ~w10312;
	assign w10449 = w50852 ^ w50868;
	assign w10345 = ~w10449;
	assign w10374 = w10345 ^ w45810;
	assign w10273 = w45956 ^ w45205;
	assign w9928 = w9958 ^ w9921;
	assign w10004 = w9925 ^ w9928;
	assign w9982 = w10004 & w10045;
	assign w9991 = w10004 & w10036;
	assign w9969 = w9987 ^ w9991;
	assign w9947 = ~w9969;
	assign w9951 = w9947 ^ w9952;
	assign w9948 = w9993 ^ w9982;
	assign w9944 = ~w9948;
	assign w10051 = w9950 ^ w9951;
	assign w45206 = ~w10051;
	assign w10504 = w45206 ^ w45810;
	assign w10235 = w45206 ^ w45877;
	assign w10510 = w10234 ^ w10235;
	assign w10416 = w45206 ^ w10238;
	assign w9997 = w10011 & w46324;
	assign w9939 = w9997 ^ w9970;
	assign w50850 = w9938 ^ w9939;
	assign w10191 = w10449 ^ w50850;
	assign w43806 = w9997 ^ w9999;
	assign w9955 = w43806 ^ w9952;
	assign w10052 = w9954 ^ w9955;
	assign w45207 = ~w10052;
	assign w10505 = w45207 ^ w45811;
	assign w10231 = w42421 ^ w45207;
	assign w9946 = w9947 ^ w9985;
	assign w9942 = w9946 ^ w43806;
	assign w9945 = w9984 ^ w9942;
	assign w10049 = w9944 ^ w9945;
	assign w9941 = w9965 ^ w9942;
	assign w50849 = w9940 ^ w9941;
	assign w10484 = w50849 ^ w50864;
	assign w10346 = ~w10484;
	assign w10343 = w10496 ^ w10346;
	assign w45211 = ~w10049;
	assign w10293 = w10486 ^ w45211;
	assign w50540 = w9900 ^ w9884;
	assign w46336 = w50540 ^ w595;
	assign w42598 = w46336 ^ w46334;
	assign w42684 = w46336 ^ w46333;
	assign w42680 = w42684 ^ w42612;
	assign w42676 = w42595 ^ w42684;
	assign w42675 = w46340 ^ w42676;
	assign w42686 = w46338 ^ w46336;
	assign w42671 = w42596 ^ w42686;
	assign w42558 = w42598 ^ w42596;
	assign w42674 = w42595 ^ w42558;
	assign w42557 = w42598 ^ w46335;
	assign w42681 = w46340 ^ w42557;
	assign w42669 = w42676 & w42680;
	assign w42601 = w42669 ^ w42598;
	assign w42668 = w42677 & w42675;
	assign w42667 = w46340 & w42681;
	assign w42663 = w42684 & w42673;
	assign w42599 = w42663 ^ w42597;
	assign w42605 = w42601 ^ w42599;
	assign w42610 = w46333 ^ w42605;
	assign w42662 = w42686 & w42671;
	assign w42619 = w42662 ^ w42668;
	assign w42660 = w42619 ^ w42610;
	assign w42571 = w42662 ^ w42663;
	assign w42618 = w42571 ^ w42572;
	assign w42617 = w42618 ^ w42600;
	assign w42659 = w42665 ^ w42617;
	assign w42661 = w42683 & w42674;
	assign w42656 = w42660 & w42659;
	assign w45155 = w42661 ^ w42664;
	assign w42574 = w42600 ^ w45155;
	assign w42658 = w42574 ^ w42599;
	assign w42655 = w42656 ^ w42658;
	assign w42614 = w42662 ^ w45155;
	assign w42570 = w42665 ^ w42614;
	assign w42652 = w46339 ^ w42570;
	assign w45158 = w42661 ^ w42667;
	assign w42573 = w42605 ^ w45158;
	assign w42616 = w46335 ^ w42573;
	assign w42651 = w42656 ^ w42616;
	assign w42650 = w42651 & w42652;
	assign w42648 = w42656 ^ w42650;
	assign w42569 = w42650 ^ w42614;
	assign w42568 = w42650 ^ w42667;
	assign w42563 = w42568 ^ w42664;
	assign w42647 = w42658 & w42648;
	assign w42645 = w42647 ^ w42655;
	assign w45157 = w42647 ^ w42665;
	assign w42639 = w45157 ^ w42617;
	assign w42628 = w42639 & w42680;
	assign w42637 = w42639 & w42676;
	assign w42606 = w46339 ^ w45157;
	assign w42646 = w42606 ^ w42569;
	assign w42636 = w42646 & w42675;
	assign w42627 = w42646 & w42677;
	assign w42649 = w42650 ^ w42658;
	assign w42635 = w42649 & w46340;
	assign w42626 = w42649 & w42681;
	assign w42611 = w45158 ^ w42596;
	assign w42657 = w42619 ^ w42611;
	assign w42654 = w42655 & w42657;
	assign w42653 = w42654 ^ w42616;
	assign w42565 = w42654 ^ w42666;
	assign w42561 = w42565 ^ w42601;
	assign w42564 = w46333 ^ w42561;
	assign w42641 = w42563 ^ w42564;
	assign w42562 = w42654 ^ w42610;
	assign w42560 = w46335 ^ w42561;
	assign w42644 = w42653 & w42645;
	assign w42609 = w42644 ^ w42619;
	assign w42643 = w42609 ^ w42611;
	assign w42567 = w42644 ^ w42668;
	assign w42559 = w42606 ^ w42567;
	assign w42566 = w42596 ^ w42559;
	assign w42642 = w42563 ^ w42566;
	assign w42640 = w42609 ^ w42562;
	assign w42638 = w42559 ^ w42560;
	assign w42634 = w42640 & w42670;
	assign w42633 = w42643 & w42682;
	assign w42632 = w42653 & w42672;
	assign w42576 = w42632 ^ w42633;
	assign w42631 = w42641 & w42673;
	assign w42630 = w42638 & w42671;
	assign w42591 = w42630 ^ w42633;
	assign w42588 = ~w42591;
	assign w42587 = w42630 ^ w42631;
	assign w42629 = w42642 & w42674;
	assign w42625 = w42640 & w42685;
	assign w42607 = w42625 ^ w42629;
	assign w42592 = w42634 ^ w42625;
	assign w42585 = ~w42607;
	assign w42624 = w42643 & w42678;
	assign w42594 = w42632 ^ w42624;
	assign w42623 = w42653 & w42679;
	assign w42584 = w42585 ^ w42623;
	assign w42622 = w42641 & w42684;
	assign w42621 = w42638 & w42686;
	assign w42620 = w42642 & w42683;
	assign w42586 = w42631 ^ w42620;
	assign w42582 = ~w42586;
	assign w45156 = w42621 ^ w42622;
	assign w42603 = w42627 ^ w45156;
	assign w42604 = w42628 ^ w42603;
	assign w42608 = w42636 ^ w42604;
	assign w42577 = w42635 ^ w42608;
	assign w50879 = w42576 ^ w42577;
	assign w10464 = w50879 ^ w50883;
	assign w10210 = w50879 ^ w10198;
	assign w42613 = w42637 ^ w42608;
	assign w42688 = w42613 ^ w42587;
	assign w42590 = w42594 ^ w45156;
	assign w42589 = w42585 ^ w42590;
	assign w42689 = w42588 ^ w42589;
	assign w45159 = w42633 ^ w42634;
	assign w50880 = w45159 ^ w42613;
	assign w10459 = w50880 ^ w50884;
	assign w10308 = ~w50880;
	assign w10323 = w10308 ^ w50876;
	assign w42615 = w42630 ^ w45159;
	assign w42581 = w42626 ^ w42615;
	assign w42578 = ~w42581;
	assign w42575 = w42631 ^ w42615;
	assign w50881 = w42604 ^ w42575;
	assign w45160 = w42635 ^ w42637;
	assign w42593 = w45160 ^ w42590;
	assign w42690 = w42592 ^ w42593;
	assign w42580 = w42584 ^ w45160;
	assign w42583 = w42622 ^ w42580;
	assign w42687 = w42582 ^ w42583;
	assign w42579 = w42603 ^ w42580;
	assign w50878 = w42578 ^ w42579;
	assign w10208 = w50878 ^ w50874;
	assign w10446 = w50877 ^ w50881;
	assign w10207 = w10446 ^ w50883;
	assign w10205 = w10446 ^ w45806;
	assign w10211 = ~w10446;
	assign w10209 = w10211 ^ w50884;
	assign w10521 = w10207 ^ w10208;
	assign w10520 = w10209 ^ w10210;
	assign w10469 = w50878 ^ w50882;
	assign w10352 = w10469 ^ w45806;
	assign w10438 = w50881 ^ w50885;
	assign w10307 = w10438 ^ w10308;
	assign w10329 = w10438 ^ w45839;
	assign w10314 = w10438 ^ w50879;
	assign w45878 = ~w42690;
	assign w10476 = w45878 ^ w45807;
	assign w10206 = w45878 ^ w45840;
	assign w10522 = w10205 ^ w10206;
	assign w45883 = ~w42687;
	assign w10454 = w45883 ^ w45812;
	assign w10350 = w10454 ^ w50884;
	assign w45884 = ~w42688;
	assign w10456 = w45839 ^ w45884;
	assign w10304 = w10456 ^ w10454;
	assign w10348 = w10456 ^ w45813;
	assign w10303 = w50881 ^ w45884;
	assign w45885 = ~w42689;
	assign w10472 = w45885 ^ w45806;
	assign w10317 = w10438 ^ w45885;
	assign w10326 = w45885 ^ w40545;
	assign w39438 = w39441 & w39439;
	assign w39349 = w39438 ^ w39450;
	assign w39437 = w39438 ^ w39400;
	assign w39428 = w39437 & w39429;
	assign w39393 = w39428 ^ w39403;
	assign w39427 = w39393 ^ w39395;
	assign w39416 = w39437 & w39456;
	assign w39417 = w39427 & w39466;
	assign w39360 = w39416 ^ w39417;
	assign w39407 = w39437 & w39463;
	assign w39351 = w39428 ^ w39452;
	assign w39343 = w39390 ^ w39351;
	assign w39350 = w39380 ^ w39343;
	assign w39426 = w39347 ^ w39350;
	assign w39413 = w39426 & w39458;
	assign w39408 = w39427 & w39462;
	assign w39378 = w39416 ^ w39408;
	assign w39345 = w39349 ^ w39385;
	assign w39348 = w46389 ^ w39345;
	assign w39425 = w39347 ^ w39348;
	assign w39415 = w39425 & w39457;
	assign w39406 = w39425 & w39468;
	assign w39404 = w39426 & w39467;
	assign w39370 = w39415 ^ w39404;
	assign w39366 = ~w39370;
	assign w39346 = w39438 ^ w39394;
	assign w39424 = w39393 ^ w39346;
	assign w39409 = w39424 & w39469;
	assign w39418 = w39424 & w39454;
	assign w39376 = w39418 ^ w39409;
	assign w45025 = w39417 ^ w39418;
	assign w39391 = w39409 ^ w39413;
	assign w39369 = ~w39391;
	assign w39368 = w39369 ^ w39407;
	assign w39364 = w39368 ^ w45026;
	assign w39344 = w46391 ^ w39345;
	assign w39422 = w39343 ^ w39344;
	assign w39414 = w39422 & w39455;
	assign w39399 = w39414 ^ w45025;
	assign w39365 = w39410 ^ w39399;
	assign w39362 = ~w39365;
	assign w39405 = w39422 & w39470;
	assign w39371 = w39414 ^ w39415;
	assign w45022 = w39405 ^ w39406;
	assign w39387 = w39411 ^ w45022;
	assign w39388 = w39412 ^ w39387;
	assign w39374 = w39378 ^ w45022;
	assign w39377 = w45026 ^ w39374;
	assign w39474 = w39376 ^ w39377;
	assign w39375 = w39414 ^ w39417;
	assign w39392 = w39420 ^ w39388;
	assign w39361 = w39419 ^ w39392;
	assign w50701 = w39360 ^ w39361;
	assign w9864 = w50697 ^ w50701;
	assign w9637 = w9639 ^ w9864;
	assign w9609 = w9612 ^ w50701;
	assign w9902 = w9609 ^ w9610;
	assign w50603 = w9902 ^ w9875;
	assign w46273 = w50603 ^ w530;
	assign w39397 = w39421 ^ w39392;
	assign w50702 = w45025 ^ w39397;
	assign w9613 = w9612 ^ w50702;
	assign w9855 = w50698 ^ w50702;
	assign w9636 = w9860 ^ w9855;
	assign w50613 = w45841 ^ w9636;
	assign w46263 = w50613 ^ w540;
	assign w9665 = w9642 ^ w9855;
	assign w50596 = w9665 ^ w9666;
	assign w39472 = w39397 ^ w39371;
	assign w46280 = w50596 ^ w523;
	assign w39372 = ~w39375;
	assign w9667 = w9658 ^ w9864;
	assign w50595 = w9667 ^ w9668;
	assign w46281 = w50595 ^ w522;
	assign w39359 = w39415 ^ w39399;
	assign w50703 = w39388 ^ w39359;
	assign w9832 = w50688 ^ w50703;
	assign w9605 = w9832 ^ w50701;
	assign w9904 = w9605 ^ w9606;
	assign w9649 = w45895 ^ w50703;
	assign w9601 = ~w9832;
	assign w9824 = w50699 ^ w50703;
	assign w9662 = w9853 ^ w9824;
	assign w50599 = w50688 ^ w9662;
	assign w9918 = ~w9824;
	assign w9641 = w9918 ^ w50697;
	assign w46277 = w50599 ^ w526;
	assign w9638 = w9918 ^ w50698;
	assign w50607 = w9649 ^ w9650;
	assign w46269 = w50607 ^ w534;
	assign w40674 = w46280 ^ w46277;
	assign w50612 = w9637 ^ w9638;
	assign w46264 = w50612 ^ w539;
	assign w9901 = w9613 ^ w9614;
	assign w50604 = w9901 ^ w9867;
	assign w46272 = w50604 ^ w531;
	assign w39363 = w39387 ^ w39364;
	assign w9646 = w9918 ^ w45835;
	assign w50700 = w39362 ^ w39363;
	assign w9656 = w9658 ^ w50700;
	assign w9602 = w9601 ^ w50700;
	assign w9905 = w9602 ^ w9603;
	assign w50587 = w9905 ^ w9864;
	assign w9874 = w50696 ^ w50700;
	assign w9640 = w9642 ^ w9874;
	assign w9687 = ~w9874;
	assign w9669 = w9889 ^ w9874;
	assign w50594 = w50685 ^ w9669;
	assign w46282 = w50594 ^ w521;
	assign w40673 = w46277 ^ w46282;
	assign w40562 = w46281 ^ w46282;
	assign w46289 = w50587 ^ w514;
	assign w50611 = w9640 ^ w9641;
	assign w46265 = w50611 ^ w538;
	assign w50602 = w9656 ^ w9657;
	assign w46274 = w50602 ^ w529;
	assign w41343 = w46269 ^ w46274;
	assign w41346 = w46274 ^ w46272;
	assign w41232 = w46273 ^ w46274;
	assign w39373 = w39369 ^ w39374;
	assign w45814 = ~w39472;
	assign w9674 = w9824 ^ w45814;
	assign w50591 = w9674 ^ w9675;
	assign w46285 = w50591 ^ w518;
	assign w9653 = w9853 ^ w45814;
	assign w9838 = w45834 ^ w45814;
	assign w9663 = w9860 ^ w9838;
	assign w9634 = w9838 ^ w9827;
	assign w50598 = w45830 ^ w9663;
	assign w46278 = w50598 ^ w525;
	assign w40588 = w46280 ^ w46278;
	assign w50615 = w50699 ^ w9634;
	assign w46261 = w50615 ^ w542;
	assign w39870 = w46264 ^ w46261;
	assign w39782 = w46263 ^ w46261;
	assign w45816 = ~w39474;
	assign w9886 = w45836 ^ w45816;
	assign w9688 = w9886 ^ w9832;
	assign w9673 = w9886 ^ w9827;
	assign w50592 = w45832 ^ w9673;
	assign w46284 = w50592 ^ w519;
	assign w40592 = w46284 ^ w46278;
	assign w50584 = w45214 ^ w9688;
	assign w9599 = w9601 ^ w45816;
	assign w9906 = w9599 ^ w9600;
	assign w9647 = w9889 ^ w9886;
	assign w9645 = ~w9647;
	assign w50609 = w9645 ^ w9646;
	assign w46267 = w50609 ^ w536;
	assign w39781 = w46267 ^ w46265;
	assign w39862 = w39781 ^ w39870;
	assign w46292 = w50584 ^ w511;
	assign w39871 = w46261 ^ w46267;
	assign w9651 = ~w9653;
	assign w50606 = w9651 ^ w9652;
	assign w46270 = w50606 ^ w533;
	assign w41258 = w46272 ^ w46270;
	assign w41344 = w46272 ^ w46269;
	assign w39473 = w39372 ^ w39373;
	assign w45815 = ~w39473;
	assign w9685 = w9687 ^ w45815;
	assign w50586 = w9685 ^ w9686;
	assign w9607 = w9831 ^ w45815;
	assign w9903 = w9607 ^ w9608;
	assign w50601 = w9903 ^ w9889;
	assign w46275 = w50601 ^ w528;
	assign w41255 = w46275 ^ w46273;
	assign w41257 = w46274 ^ w41255;
	assign w41345 = w46269 ^ w46275;
	assign w41336 = w41255 ^ w41344;
	assign w41272 = w46275 ^ w46274;
	assign w46290 = w50586 ^ w513;
	assign w42549 = w46285 ^ w46290;
	assign w41333 = w46270 ^ w41257;
	assign w41323 = w41344 & w41333;
	assign w41259 = w41323 ^ w41257;
	assign w9878 = w45835 ^ w45815;
	assign w9671 = w9890 ^ w9878;
	assign w50585 = w9906 ^ w9878;
	assign w9643 = w9882 ^ w9878;
	assign w46291 = w50585 ^ w512;
	assign w42551 = w46285 ^ w46291;
	assign w42461 = w46291 ^ w46289;
	assign w9670 = w9671 ^ w9672;
	assign w42463 = w46290 ^ w42461;
	assign w50610 = w50696 ^ w9643;
	assign w50593 = ~w9670;
	assign w46283 = w50593 ^ w520;
	assign w40585 = w46283 ^ w46281;
	assign w40587 = w46282 ^ w40585;
	assign w40663 = w46278 ^ w40587;
	assign w40653 = w40674 & w40663;
	assign w40666 = w40585 ^ w40674;
	assign w40602 = w46283 ^ w46282;
	assign w40665 = w46284 ^ w40666;
	assign w40670 = w40674 ^ w40602;
	assign w40659 = w40666 & w40670;
	assign w40589 = w40653 ^ w40587;
	assign w46266 = w50610 ^ w537;
	assign w39798 = w46267 ^ w46266;
	assign w39866 = w39870 ^ w39798;
	assign w39872 = w46266 ^ w46264;
	assign w39783 = w46266 ^ w39781;
	assign w39856 = w46263 ^ w39783;
	assign w39852 = w39871 & w39856;
	assign w39786 = w39852 ^ w39782;
	assign w39758 = w46265 ^ w46266;
	assign w39855 = w39862 & w39866;
	assign w40591 = w40659 ^ w40588;
	assign w39869 = w46261 ^ w46266;
	assign w39857 = w39782 ^ w39872;
	assign w39848 = w39872 & w39857;
	assign w42478 = w46291 ^ w46290;
	assign w40595 = w40591 ^ w40589;
	assign w40600 = w46277 ^ w40595;
	assign w40675 = w46277 ^ w46283;
	assign w42438 = w46289 ^ w46290;
	assign w41340 = w41344 ^ w41272;
	assign w41329 = w41336 & w41340;
	assign w41261 = w41329 ^ w41258;
	assign w40662 = w40592 ^ w40587;
	assign w39367 = w39406 ^ w39364;
	assign w39471 = w39366 ^ w39367;
	assign w45821 = ~w39471;
	assign w9849 = w45841 ^ w45821;
	assign w9684 = w9849 ^ w50702;
	assign w9682 = ~w9684;
	assign w9664 = w9867 ^ w9849;
	assign w9654 = w9860 ^ w45821;
	assign w50605 = w9654 ^ w9655;
	assign w9677 = w9838 ^ w45821;
	assign w9676 = w9677 ^ w9678;
	assign w50590 = ~w9676;
	assign w46286 = w50590 ^ w517;
	assign w46271 = w50605 ^ w532;
	assign w50589 = w9682 ^ w9683;
	assign w46287 = w50589 ^ w516;
	assign w42462 = w46287 ^ w46285;
	assign w42536 = w46287 ^ w42463;
	assign w9635 = w9853 ^ w9849;
	assign w41330 = w46271 ^ w41257;
	assign w41326 = w41345 & w41330;
	assign w41256 = w46271 ^ w46269;
	assign w41331 = w41256 ^ w41346;
	assign w41322 = w41346 & w41331;
	assign w41231 = w41322 ^ w41323;
	assign w41278 = w41231 ^ w41232;
	assign w41260 = w41326 ^ w41256;
	assign w41277 = w41278 ^ w41260;
	assign w42539 = w46286 ^ w42463;
	assign w41217 = w41258 ^ w46271;
	assign w42532 = w42551 & w42536;
	assign w42466 = w42532 ^ w42462;
	assign w41218 = w41258 ^ w41256;
	assign w42468 = w46292 ^ w46286;
	assign w42538 = w42468 ^ w42463;
	assign w42548 = w46287 ^ w42468;
	assign w42545 = w42462 ^ w42468;
	assign w42530 = w42545 & w42538;
	assign w42543 = w42478 ^ w42545;
	assign w41334 = w41255 ^ w41218;
	assign w41321 = w41343 & w41334;
	assign w50597 = w45837 ^ w9664;
	assign w46279 = w50597 ^ w524;
	assign w40547 = w40588 ^ w46279;
	assign w40660 = w46279 ^ w40587;
	assign w40586 = w46279 ^ w46277;
	assign w40548 = w40588 ^ w40586;
	assign w40664 = w40585 ^ w40548;
	assign w40651 = w40673 & w40664;
	assign w40669 = w40586 ^ w40592;
	assign w40667 = w40602 ^ w40669;
	assign w40654 = w40669 & w40662;
	assign w40658 = w40667 & w40665;
	assign w40656 = w40675 & w40660;
	assign w45073 = w40651 ^ w40654;
	assign w40672 = w46279 ^ w40592;
	assign w40668 = w46283 ^ w40672;
	assign w40590 = w40656 ^ w40586;
	assign w40564 = w40590 ^ w45073;
	assign w40648 = w40564 ^ w40589;
	assign w40655 = w40672 & w40668;
	assign w40671 = w46284 ^ w40547;
	assign w40657 = w46284 & w40671;
	assign w45072 = w40651 ^ w40657;
	assign w40601 = w45072 ^ w40586;
	assign w40563 = w40595 ^ w45072;
	assign w40606 = w46279 ^ w40563;
	assign w42544 = w46291 ^ w42548;
	assign w42531 = w42548 & w42544;
	assign w40676 = w46282 ^ w46280;
	assign w40661 = w40586 ^ w40676;
	assign w40652 = w40676 & w40661;
	assign w40561 = w40652 ^ w40653;
	assign w40608 = w40561 ^ w40562;
	assign w40607 = w40608 ^ w40590;
	assign w40604 = w40652 ^ w45073;
	assign w40560 = w40655 ^ w40604;
	assign w40642 = w46283 ^ w40560;
	assign w40649 = w40655 ^ w40607;
	assign w40609 = w40652 ^ w40658;
	assign w40650 = w40609 ^ w40600;
	assign w40646 = w40650 & w40649;
	assign w40641 = w40646 ^ w40606;
	assign w40640 = w40641 & w40642;
	assign w40638 = w40646 ^ w40640;
	assign w40558 = w40640 ^ w40657;
	assign w40553 = w40558 ^ w40654;
	assign w40637 = w40648 & w40638;
	assign w40639 = w40640 ^ w40648;
	assign w40616 = w40639 & w40671;
	assign w45076 = w40637 ^ w40655;
	assign w40629 = w45076 ^ w40607;
	assign w40627 = w40629 & w40666;
	assign w40618 = w40629 & w40670;
	assign w40596 = w46283 ^ w45076;
	assign w40625 = w40639 & w46284;
	assign w45075 = w40625 ^ w40627;
	assign w40645 = w40646 ^ w40648;
	assign w40635 = w40637 ^ w40645;
	assign w40647 = w40609 ^ w40601;
	assign w40644 = w40647 & w40645;
	assign w40552 = w40644 ^ w40600;
	assign w40643 = w40644 ^ w40606;
	assign w40622 = w40643 & w40662;
	assign w40613 = w40643 & w40669;
	assign w40555 = w40644 ^ w40656;
	assign w40551 = w40555 ^ w40591;
	assign w40554 = w46277 ^ w40551;
	assign w40631 = w40553 ^ w40554;
	assign w40550 = w46279 ^ w40551;
	assign w40634 = w40643 & w40635;
	assign w40557 = w40634 ^ w40658;
	assign w40549 = w40596 ^ w40557;
	assign w40556 = w40586 ^ w40549;
	assign w40632 = w40553 ^ w40556;
	assign w40610 = w40632 & w40673;
	assign w40619 = w40632 & w40664;
	assign w40628 = w40549 ^ w40550;
	assign w40611 = w40628 & w40676;
	assign w40620 = w40628 & w40661;
	assign w40612 = w40631 & w40674;
	assign w43611 = w40611 ^ w40612;
	assign w40599 = w40634 ^ w40609;
	assign w40630 = w40599 ^ w40552;
	assign w40615 = w40630 & w40675;
	assign w40624 = w40630 & w40660;
	assign w40633 = w40599 ^ w40601;
	assign w40614 = w40633 & w40668;
	assign w40584 = w40622 ^ w40614;
	assign w40623 = w40633 & w40672;
	assign w40581 = w40620 ^ w40623;
	assign w40578 = ~w40581;
	assign w40566 = w40622 ^ w40623;
	assign w40580 = w40584 ^ w43611;
	assign w40583 = w45075 ^ w40580;
	assign w45074 = w40623 ^ w40624;
	assign w40582 = w40624 ^ w40615;
	assign w40680 = w40582 ^ w40583;
	assign w40597 = w40615 ^ w40619;
	assign w40575 = ~w40597;
	assign w40574 = w40575 ^ w40613;
	assign w40570 = w40574 ^ w45075;
	assign w40573 = w40612 ^ w40570;
	assign w40579 = w40575 ^ w40580;
	assign w40679 = w40578 ^ w40579;
	assign w40621 = w40631 & w40663;
	assign w40577 = w40620 ^ w40621;
	assign w40576 = w40621 ^ w40610;
	assign w40572 = ~w40576;
	assign w40677 = w40572 ^ w40573;
	assign w10311 = w50866 ^ w40677;
	assign w50726 = w10310 ^ w10311;
	assign w46223 = w50726 ^ w708;
	assign w10369 = w45875 ^ w40677;
	assign w50856 = ~w40677;
	assign w10494 = w45211 ^ w50856;
	assign w10358 = w10494 ^ w10493;
	assign w10384 = w10494 ^ w10486;
	assign w50735 = w45205 ^ w10384;
	assign w46214 = w50735 ^ w717;
	assign w10370 = w10494 ^ w45817;
	assign w50750 = w45875 ^ w10358;
	assign w46199 = w50750 ^ w732;
	assign w45844 = ~w40679;
	assign w10483 = w45844 ^ w50859;
	assign w50746 = w10510 ^ w10483;
	assign w10378 = w10484 ^ w10483;
	assign w10415 = w10346 ^ w45844;
	assign w50731 = w10415 ^ w10416;
	assign w46218 = w50731 ^ w713;
	assign w46203 = w50746 ^ w728;
	assign w10373 = w10505 ^ w10483;
	assign w10372 = w10373 ^ w10374;
	assign w50722 = ~w10372;
	assign w46227 = w50722 ^ w704;
	assign w45845 = ~w40680;
	assign w10482 = w45845 ^ w45877;
	assign w10365 = w10482 ^ w10441;
	assign w50745 = w45207 ^ w10365;
	assign w46204 = w50745 ^ w727;
	assign w10434 = w10482 ^ w10449;
	assign w50721 = w45811 ^ w10434;
	assign w46228 = w50721 ^ w703;
	assign w40605 = w40620 ^ w45074;
	assign w40565 = w40621 ^ w40605;
	assign w40571 = w40616 ^ w40605;
	assign w40568 = ~w40571;
	assign w40559 = w40640 ^ w40604;
	assign w40636 = w40596 ^ w40559;
	assign w40626 = w40636 & w40665;
	assign w40617 = w40636 & w40667;
	assign w40593 = w40617 ^ w43611;
	assign w40569 = w40593 ^ w40570;
	assign w50853 = w40568 ^ w40569;
	assign w10481 = w50853 ^ w50860;
	assign w10357 = w10504 ^ w10481;
	assign w40594 = w40618 ^ w40593;
	assign w40598 = w40626 ^ w40594;
	assign w40603 = w40627 ^ w40598;
	assign w50855 = w45074 ^ w40603;
	assign w10371 = w50862 ^ w50855;
	assign w40678 = w40603 ^ w40577;
	assign w10367 = w45876 ^ w40678;
	assign w10294 = w45817 ^ w40678;
	assign w50858 = w40594 ^ w40565;
	assign w10274 = w39338 ^ w50858;
	assign w50728 = w10273 ^ w10274;
	assign w46221 = w50728 ^ w710;
	assign w2177 = w46221 ^ w46227;
	assign w10442 = w50852 ^ w50858;
	assign w10232 = w10442 ^ w50850;
	assign w10257 = w10505 ^ w10442;
	assign w50729 = w45877 ^ w10257;
	assign w10355 = w10486 ^ w10442;
	assign w46220 = w50729 ^ w711;
	assign w50752 = w50863 ^ w10355;
	assign w46197 = w50752 ^ w734;
	assign w2579 = w46197 ^ w46203;
	assign w2072 = w46223 ^ w46221;
	assign w10497 = w50851 ^ w50855;
	assign w10385 = w10497 ^ w10489;
	assign w10361 = w10497 ^ w10496;
	assign w10359 = ~w10361;
	assign w50749 = w10359 ^ w10360;
	assign w46200 = w50749 ^ w731;
	assign w10192 = w50865 ^ w50855;
	assign w2228 = w46220 ^ w46214;
	assign w2490 = w46199 ^ w46197;
	assign w50742 = w10370 ^ w10371;
	assign w10443 = w50858 ^ w50863;
	assign w10377 = ~w10443;
	assign w10376 = w10377 ^ w50865;
	assign w10381 = w10377 ^ w45844;
	assign w10228 = w10443 ^ w50866;
	assign w50734 = w45211 ^ w10385;
	assign w46215 = w50734 ^ w716;
	assign w2308 = w46215 ^ w2228;
	assign w50723 = w50864 ^ w10357;
	assign w46226 = w50723 ^ w705;
	assign w2175 = w46221 ^ w46226;
	assign w2055 = w46227 ^ w46226;
	assign w50857 = ~w40678;
	assign w10492 = w45205 ^ w50857;
	assign w10383 = w10492 ^ w10441;
	assign w10368 = w10492 ^ w39338;
	assign w50743 = w10368 ^ w10369;
	assign w46206 = w50743 ^ w725;
	assign w40567 = w40625 ^ w40598;
	assign w50854 = w40566 ^ w40567;
	assign w10506 = w50850 ^ w50854;
	assign w50748 = w10509 ^ w10506;
	assign w46201 = w50748 ^ w730;
	assign w2489 = w46203 ^ w46201;
	assign w10344 = w10345 ^ w50854;
	assign w10388 = ~w10506;
	assign w10386 = w10388 ^ w10493;
	assign w10229 = w50861 ^ w50854;
	assign w10513 = w10228 ^ w10229;
	assign w10364 = ~w10481;
	assign w10362 = w10364 ^ w50849;
	assign w50747 = w10362 ^ w10363;
	assign w46202 = w50747 ^ w729;
	assign w2506 = w46203 ^ w46202;
	assign w2577 = w46197 ^ w46202;
	assign w2580 = w46202 ^ w46200;
	assign w2565 = w2490 ^ w2580;
	assign w2556 = w2580 & w2565;
	assign w2466 = w46201 ^ w46202;
	assign w10375 = w10506 ^ w10364;
	assign w2491 = w46202 ^ w2489;
	assign w2564 = w46199 ^ w2491;
	assign w2560 = w2579 & w2564;
	assign w10233 = w50849 ^ w50853;
	assign w10511 = w10232 ^ w10233;
	assign w50732 = w10511 ^ w10496;
	assign w46217 = w50732 ^ w714;
	assign w2198 = w46217 ^ w46218;
	assign w50736 = w50852 ^ w10383;
	assign w46213 = w50736 ^ w718;
	assign w2222 = w46215 ^ w46213;
	assign w2305 = w2222 ^ w2228;
	assign w2309 = w46213 ^ w46218;
	assign w50740 = w10375 ^ w10376;
	assign w46209 = w50740 ^ w722;
	assign w50724 = w10343 ^ w10344;
	assign w46225 = w50724 ^ w706;
	assign w2096 = w46225 ^ w46226;
	assign w2073 = w46227 ^ w46225;
	assign w2071 = w46226 ^ w2073;
	assign w2162 = w46223 ^ w2071;
	assign w2158 = w2177 & w2162;
	assign w2068 = w2158 ^ w2072;
	assign w2494 = w2560 ^ w2490;
	assign w10382 = w10505 ^ w10443;
	assign w50737 = w45845 ^ w10382;
	assign w46212 = w50737 ^ w719;
	assign w2362 = w46212 ^ w46206;
	assign w50739 = w50853 ^ w10378;
	assign w46210 = w50739 ^ w721;
	assign w2332 = w46209 ^ w46210;
	assign w10528 = w10191 ^ w10192;
	assign w10292 = w10293 ^ w10294;
	assign w50727 = ~w10292;
	assign w46222 = w50727 ^ w709;
	assign w2165 = w46222 ^ w2071;
	assign w2066 = w46228 ^ w46222;
	assign w2164 = w2066 ^ w2071;
	assign w2174 = w46223 ^ w2066;
	assign w2170 = w46227 ^ w2174;
	assign w2171 = w2072 ^ w2066;
	assign w2169 = w2055 ^ w2171;
	assign w2156 = w2171 & w2164;
	assign w2157 = w2174 & w2170;
	assign w50725 = w10528 ^ w10493;
	assign w46224 = w50725 ^ w707;
	assign w2178 = w46226 ^ w46224;
	assign w2163 = w2072 ^ w2178;
	assign w2154 = w2178 & w2163;
	assign w2070 = w46224 ^ w46222;
	assign w2110 = w2070 ^ w2072;
	assign w2166 = w2073 ^ w2110;
	assign w2153 = w2175 & w2166;
	assign w43620 = w2153 ^ w2156;
	assign w2053 = w2154 ^ w43620;
	assign w2098 = w2157 ^ w2053;
	assign w2094 = w2068 ^ w43620;
	assign w2111 = w2070 ^ w46223;
	assign w2173 = w46228 ^ w2111;
	assign w2159 = w46228 & w2173;
	assign w43619 = w2153 ^ w2159;
	assign w2056 = w43619 ^ w2072;
	assign w2144 = w46227 ^ w2098;
	assign w2176 = w46224 ^ w46221;
	assign w2168 = w2073 ^ w2176;
	assign w2167 = w46228 ^ w2168;
	assign w2160 = w2169 & w2167;
	assign w2155 = w2176 & w2165;
	assign w2062 = w2154 ^ w2160;
	assign w2149 = w2062 ^ w2056;
	assign w2069 = w2155 ^ w2071;
	assign w2150 = w2094 ^ w2069;
	assign w2578 = w46200 ^ w46197;
	assign w2574 = w2578 ^ w2506;
	assign w2172 = w2176 ^ w2055;
	assign w2161 = w2168 & w2172;
	assign w2067 = w2161 ^ w2070;
	assign w2063 = w2067 ^ w2069;
	assign w2057 = w46221 ^ w2063;
	assign w2095 = w2063 ^ w43619;
	assign w2051 = w46223 ^ w2095;
	assign w2152 = w2062 ^ w2057;
	assign w2570 = w2489 ^ w2578;
	assign w2563 = w2570 & w2574;
	assign w2569 = w46204 ^ w2570;
	assign w50741 = w10513 ^ w10497;
	assign w46208 = w50741 ^ w723;
	assign w2358 = w46208 ^ w46206;
	assign w2446 = w46210 ^ w46208;
	assign w10356 = w10492 ^ w10489;
	assign w50751 = w45876 ^ w10356;
	assign w46198 = w50751 ^ w733;
	assign w2567 = w46198 ^ w2491;
	assign w2557 = w2578 & w2567;
	assign w2493 = w2557 ^ w2491;
	assign w2496 = w46204 ^ w46198;
	assign w2576 = w46199 ^ w2496;
	assign w2573 = w2490 ^ w2496;
	assign w2571 = w2506 ^ w2573;
	assign w2572 = w46203 ^ w2576;
	assign w2559 = w2576 & w2572;
	assign w2562 = w2571 & w2569;
	assign w2513 = w2556 ^ w2562;
	assign w2492 = w46200 ^ w46198;
	assign w2495 = w2563 ^ w2492;
	assign w2499 = w2495 ^ w2493;
	assign w2504 = w46197 ^ w2499;
	assign w2554 = w2513 ^ w2504;
	assign w2451 = w2492 ^ w46199;
	assign w2575 = w46204 ^ w2451;
	assign w2561 = w46204 & w2575;
	assign w2566 = w2496 ^ w2491;
	assign w2558 = w2573 & w2566;
	assign w2465 = w2556 ^ w2557;
	assign w2512 = w2465 ^ w2466;
	assign w2511 = w2512 ^ w2494;
	assign w2553 = w2559 ^ w2511;
	assign w2550 = w2554 & w2553;
	assign w2452 = w2492 ^ w2490;
	assign w2568 = w2489 ^ w2452;
	assign w2555 = w2577 & w2568;
	assign w43637 = w2555 ^ w2558;
	assign w43636 = w2555 ^ w2561;
	assign w2467 = w2499 ^ w43636;
	assign w2505 = w43636 ^ w2490;
	assign w2551 = w2513 ^ w2505;
	assign w2508 = w2556 ^ w43637;
	assign w2510 = w46199 ^ w2467;
	assign w2545 = w2550 ^ w2510;
	assign w2464 = w2559 ^ w2508;
	assign w2546 = w46203 ^ w2464;
	assign w2544 = w2545 & w2546;
	assign w2463 = w2544 ^ w2508;
	assign w2542 = w2550 ^ w2544;
	assign w2462 = w2544 ^ w2561;
	assign w2457 = w2462 ^ w2558;
	assign w2097 = w2154 ^ w2155;
	assign w2049 = w2097 ^ w2096;
	assign w2050 = w2049 ^ w2068;
	assign w2151 = w2157 ^ w2050;
	assign w2148 = w2152 & w2151;
	assign w2147 = w2148 ^ w2150;
	assign w2143 = w2148 ^ w2051;
	assign w2146 = w2147 & w2149;
	assign w2103 = w2146 ^ w2158;
	assign w2107 = w2103 ^ w2067;
	assign w2106 = w2146 ^ w2057;
	assign w2108 = w46223 ^ w2107;
	assign w2104 = w46221 ^ w2107;
	assign w2142 = w2143 & w2144;
	assign w2100 = w2142 ^ w2159;
	assign w2105 = w2100 ^ w2156;
	assign w2133 = w2105 ^ w2104;
	assign w2123 = w2133 & w2165;
	assign w2140 = w2148 ^ w2142;
	assign w2139 = w2150 & w2140;
	assign w2137 = w2139 ^ w2147;
	assign w2141 = w2142 ^ w2150;
	assign w2099 = w2142 ^ w2053;
	assign w2118 = w2141 & w2173;
	assign w43624 = w2139 ^ w2157;
	assign w2061 = w46227 ^ w43624;
	assign w2138 = w2061 ^ w2099;
	assign w2128 = w2138 & w2167;
	assign w2119 = w2138 & w2169;
	assign w2131 = w43624 ^ w2050;
	assign w2129 = w2131 & w2168;
	assign w2114 = w2133 & w2176;
	assign w2145 = w2146 ^ w2051;
	assign w2136 = w2145 & w2137;
	assign w2101 = w2136 ^ w2160;
	assign w2115 = w2145 & w2171;
	assign w2124 = w2145 & w2164;
	assign w2109 = w2061 ^ w2101;
	assign w2130 = w2109 ^ w2108;
	assign w2113 = w2130 & w2178;
	assign w2122 = w2130 & w2163;
	assign w43621 = w2113 ^ w2114;
	assign w2065 = w2119 ^ w43621;
	assign w2102 = w2072 ^ w2109;
	assign w2134 = w2105 ^ w2102;
	assign w2112 = w2134 & w2175;
	assign w2121 = w2134 & w2166;
	assign w2082 = w2123 ^ w2112;
	assign w2086 = ~w2082;
	assign w2081 = w2122 ^ w2123;
	assign w2058 = w2136 ^ w2062;
	assign w2135 = w2058 ^ w2056;
	assign w2125 = w2135 & w2174;
	assign w2092 = w2124 ^ w2125;
	assign w2116 = w2135 & w2170;
	assign w2077 = w2122 ^ w2125;
	assign w2080 = ~w2077;
	assign w2132 = w2058 ^ w2106;
	assign w2126 = w2132 & w2162;
	assign w43622 = w2125 ^ w2126;
	assign w2052 = w2122 ^ w43622;
	assign w2093 = w2123 ^ w2052;
	assign w2087 = w2118 ^ w2052;
	assign w2090 = ~w2087;
	assign w2074 = w2124 ^ w2116;
	assign w2078 = w2074 ^ w43621;
	assign w2117 = w2132 & w2177;
	assign w2076 = w2126 ^ w2117;
	assign w2060 = w2117 ^ w2121;
	assign w2083 = ~w2060;
	assign w2079 = w2083 ^ w2078;
	assign w2181 = w2080 ^ w2079;
	assign w46070 = ~w2181;
	assign w51019 = w46070 ^ w736;
	assign w2084 = w2083 ^ w2115;
	assign w46207 = w50742 ^ w724;
	assign w2442 = w46207 ^ w2362;
	assign w2317 = w2358 ^ w46207;
	assign w2441 = w46212 ^ w2317;
	assign w2427 = w46212 & w2441;
	assign w2468 = w2494 ^ w43637;
	assign w2552 = w2468 ^ w2493;
	assign w2549 = w2550 ^ w2552;
	assign w2541 = w2552 & w2542;
	assign w2548 = w2551 & w2549;
	assign w2456 = w2548 ^ w2504;
	assign w2543 = w2544 ^ w2552;
	assign w2520 = w2543 & w2575;
	assign w2529 = w2543 & w46204;
	assign w2539 = w2541 ^ w2549;
	assign w2547 = w2548 ^ w2510;
	assign w2517 = w2547 & w2573;
	assign w2538 = w2547 & w2539;
	assign w2503 = w2538 ^ w2513;
	assign w2459 = w2548 ^ w2560;
	assign w2455 = w2459 ^ w2495;
	assign w2458 = w46197 ^ w2455;
	assign w2535 = w2457 ^ w2458;
	assign w2525 = w2535 & w2567;
	assign w2516 = w2535 & w2578;
	assign w2537 = w2503 ^ w2505;
	assign w2518 = w2537 & w2572;
	assign w2527 = w2537 & w2576;
	assign w2526 = w2547 & w2566;
	assign w2470 = w2526 ^ w2527;
	assign w2488 = w2526 ^ w2518;
	assign w43641 = w2541 ^ w2559;
	assign w2500 = w46203 ^ w43641;
	assign w2540 = w2500 ^ w2463;
	assign w2521 = w2540 & w2571;
	assign w2533 = w43641 ^ w2511;
	assign w2531 = w2533 & w2570;
	assign w43640 = w2529 ^ w2531;
	assign w2522 = w2533 & w2574;
	assign w2534 = w2503 ^ w2456;
	assign w2528 = w2534 & w2564;
	assign w43639 = w2527 ^ w2528;
	assign w2454 = w46199 ^ w2455;
	assign w2519 = w2534 & w2579;
	assign w2486 = w2528 ^ w2519;
	assign w2530 = w2540 & w2569;
	assign w2461 = w2538 ^ w2562;
	assign w2453 = w2500 ^ w2461;
	assign w2532 = w2453 ^ w2454;
	assign w2515 = w2532 & w2580;
	assign w2524 = w2532 & w2565;
	assign w2509 = w2524 ^ w43639;
	assign w2475 = w2520 ^ w2509;
	assign w2472 = ~w2475;
	assign w2469 = w2525 ^ w2509;
	assign w2481 = w2524 ^ w2525;
	assign w43638 = w2515 ^ w2516;
	assign w2484 = w2488 ^ w43638;
	assign w2487 = w43640 ^ w2484;
	assign w2584 = w2486 ^ w2487;
	assign w45997 = ~w2584;
	assign w50946 = w45997 ^ w855;
	assign w2460 = w2490 ^ w2453;
	assign w2536 = w2457 ^ w2460;
	assign w2485 = w2524 ^ w2527;
	assign w2482 = ~w2485;
	assign w2497 = w2521 ^ w43638;
	assign w2498 = w2522 ^ w2497;
	assign w2502 = w2530 ^ w2498;
	assign w2507 = w2531 ^ w2502;
	assign w46001 = w43639 ^ w2507;
	assign w2582 = w2507 ^ w2481;
	assign w46004 = w2498 ^ w2469;
	assign w50953 = w46004 ^ w862;
	assign w2471 = w2529 ^ w2502;
	assign w46000 = w2470 ^ w2471;
	assign w50949 = w46000 ^ w858;
	assign w2514 = w2536 & w2577;
	assign w2480 = w2525 ^ w2514;
	assign w2476 = ~w2480;
	assign w2523 = w2536 & w2568;
	assign w2501 = w2519 ^ w2523;
	assign w2479 = ~w2501;
	assign w2478 = w2479 ^ w2517;
	assign w2474 = w2478 ^ w43640;
	assign w2477 = w2516 ^ w2474;
	assign w2473 = w2497 ^ w2474;
	assign w45999 = w2472 ^ w2473;
	assign w50948 = w45999 ^ w857;
	assign w2483 = w2479 ^ w2484;
	assign w2581 = w2476 ^ w2477;
	assign w46002 = ~w2581;
	assign w2583 = w2482 ^ w2483;
	assign w45998 = ~w2583;
	assign w50947 = w45998 ^ w856;
	assign w46003 = ~w2582;
	assign w50952 = w46003 ^ w861;
	assign w50950 = w46001 ^ w859;
	assign w50951 = w46002 ^ w860;
	assign w50588 = w9904 ^ w9855;
	assign w46288 = w50588 ^ w515;
	assign w42550 = w46288 ^ w46285;
	assign w42546 = w42550 ^ w42478;
	assign w42542 = w42461 ^ w42550;
	assign w42541 = w46292 ^ w42542;
	assign w42535 = w42542 & w42546;
	assign w42529 = w42550 & w42539;
	assign w42534 = w42543 & w42541;
	assign w42464 = w46288 ^ w46286;
	assign w42424 = w42464 ^ w42462;
	assign w42540 = w42461 ^ w42424;
	assign w42527 = w42549 & w42540;
	assign w42423 = w42464 ^ w46287;
	assign w42547 = w46292 ^ w42423;
	assign w42533 = w46292 & w42547;
	assign w45150 = w42527 ^ w42533;
	assign w42477 = w45150 ^ w42462;
	assign w42465 = w42529 ^ w42463;
	assign w45151 = w42527 ^ w42530;
	assign w42467 = w42535 ^ w42464;
	assign w42471 = w42467 ^ w42465;
	assign w42439 = w42471 ^ w45150;
	assign w42482 = w46287 ^ w42439;
	assign w42440 = w42466 ^ w45151;
	assign w42476 = w46285 ^ w42471;
	assign w42552 = w46290 ^ w46288;
	assign w42537 = w42462 ^ w42552;
	assign w42528 = w42552 & w42537;
	assign w42480 = w42528 ^ w45151;
	assign w42485 = w42528 ^ w42534;
	assign w42526 = w42485 ^ w42476;
	assign w42523 = w42485 ^ w42477;
	assign w42437 = w42528 ^ w42529;
	assign w42436 = w42531 ^ w42480;
	assign w42518 = w46291 ^ w42436;
	assign w42524 = w42440 ^ w42465;
	assign w42484 = w42437 ^ w42438;
	assign w42483 = w42484 ^ w42466;
	assign w42525 = w42531 ^ w42483;
	assign w42522 = w42526 & w42525;
	assign w42517 = w42522 ^ w42482;
	assign w42516 = w42517 & w42518;
	assign w42435 = w42516 ^ w42480;
	assign w42434 = w42516 ^ w42533;
	assign w42514 = w42522 ^ w42516;
	assign w42513 = w42524 & w42514;
	assign w42515 = w42516 ^ w42524;
	assign w42501 = w42515 & w46292;
	assign w42429 = w42434 ^ w42530;
	assign w45154 = w42513 ^ w42531;
	assign w42472 = w46291 ^ w45154;
	assign w42512 = w42472 ^ w42435;
	assign w42493 = w42512 & w42543;
	assign w42505 = w45154 ^ w42483;
	assign w42494 = w42505 & w42546;
	assign w42503 = w42505 & w42542;
	assign w45153 = w42501 ^ w42503;
	assign w42502 = w42512 & w42541;
	assign w42492 = w42515 & w42547;
	assign w42521 = w42522 ^ w42524;
	assign w42511 = w42513 ^ w42521;
	assign w42520 = w42523 & w42521;
	assign w42431 = w42520 ^ w42532;
	assign w42427 = w42431 ^ w42467;
	assign w42519 = w42520 ^ w42482;
	assign w42489 = w42519 & w42545;
	assign w42510 = w42519 & w42511;
	assign w42433 = w42510 ^ w42534;
	assign w42425 = w42472 ^ w42433;
	assign w42432 = w42462 ^ w42425;
	assign w42508 = w42429 ^ w42432;
	assign w42486 = w42508 & w42549;
	assign w42495 = w42508 & w42540;
	assign w42430 = w46285 ^ w42427;
	assign w42507 = w42429 ^ w42430;
	assign w42497 = w42507 & w42539;
	assign w42452 = w42497 ^ w42486;
	assign w42448 = ~w42452;
	assign w42428 = w42520 ^ w42476;
	assign w42426 = w46287 ^ w42427;
	assign w42498 = w42519 & w42538;
	assign w42504 = w42425 ^ w42426;
	assign w42496 = w42504 & w42537;
	assign w42475 = w42510 ^ w42485;
	assign w42506 = w42475 ^ w42428;
	assign w42509 = w42475 ^ w42477;
	assign w42499 = w42509 & w42548;
	assign w42442 = w42498 ^ w42499;
	assign w42457 = w42496 ^ w42499;
	assign w42500 = w42506 & w42536;
	assign w45152 = w42499 ^ w42500;
	assign w42481 = w42496 ^ w45152;
	assign w42441 = w42497 ^ w42481;
	assign w42447 = w42492 ^ w42481;
	assign w42444 = ~w42447;
	assign w42491 = w42506 & w42551;
	assign w42473 = w42491 ^ w42495;
	assign w42458 = w42500 ^ w42491;
	assign w42490 = w42509 & w42544;
	assign w42460 = w42498 ^ w42490;
	assign w42488 = w42507 & w42550;
	assign w42487 = w42504 & w42552;
	assign w43617 = w42487 ^ w42488;
	assign w42469 = w42493 ^ w43617;
	assign w42470 = w42494 ^ w42469;
	assign w42474 = w42502 ^ w42470;
	assign w42443 = w42501 ^ w42474;
	assign w50870 = w42442 ^ w42443;
	assign w10200 = w50876 ^ w50870;
	assign w10471 = w50870 ^ w50875;
	assign w10335 = ~w10471;
	assign w10333 = w10335 ^ w10459;
	assign w42456 = w42460 ^ w43617;
	assign w50772 = w10521 ^ w10471;
	assign w46177 = w50772 ^ w690;
	assign w50872 = w42470 ^ w42441;
	assign w10439 = w50872 ^ w50877;
	assign w10319 = w10456 ^ w10439;
	assign w50776 = w50885 ^ w10319;
	assign w46173 = w50776 ^ w694;
	assign w10302 = w10439 ^ w45813;
	assign w50784 = w10302 ^ w10303;
	assign w46165 = w50784 ^ w702;
	assign w10448 = w50872 ^ w50885;
	assign w10354 = w10476 ^ w10448;
	assign w50753 = w45840 ^ w10354;
	assign w10199 = w10448 ^ w50883;
	assign w10525 = w10199 ^ w10200;
	assign w46196 = w50753 ^ w671;
	assign w50757 = w10525 ^ w10459;
	assign w46192 = w50757 ^ w675;
	assign w10342 = w10476 ^ w10439;
	assign w10313 = w10471 ^ w10469;
	assign w50780 = w10313 ^ w10314;
	assign w46169 = w50780 ^ w698;
	assign w10195 = ~w10448;
	assign w10193 = w10195 ^ w45807;
	assign w42459 = w45153 ^ w42456;
	assign w42556 = w42458 ^ w42459;
	assign w42451 = ~w42473;
	assign w42455 = w42451 ^ w42456;
	assign w42450 = w42451 ^ w42489;
	assign w42446 = w42450 ^ w45153;
	assign w42449 = w42488 ^ w42446;
	assign w42553 = w42448 ^ w42449;
	assign w42445 = w42469 ^ w42446;
	assign w50869 = w42444 ^ w42445;
	assign w10474 = w50869 ^ w50874;
	assign w10327 = ~w10474;
	assign w10336 = w10327 ^ w10464;
	assign w10325 = w10327 ^ w50882;
	assign w10315 = w10474 ^ w10472;
	assign w50779 = w50878 ^ w10315;
	assign w46170 = w50779 ^ w697;
	assign w2979 = w46165 ^ w46170;
	assign w2868 = w46169 ^ w46170;
	assign w50771 = w10325 ^ w10326;
	assign w46178 = w50771 ^ w689;
	assign w42281 = w46173 ^ w46178;
	assign w42170 = w46177 ^ w46178;
	assign w10197 = w10198 ^ w50869;
	assign w10196 = w10195 ^ w50882;
	assign w10526 = w10196 ^ w10197;
	assign w50756 = w10526 ^ w10464;
	assign w46193 = w50756 ^ w674;
	assign w42454 = ~w42457;
	assign w42555 = w42454 ^ w42455;
	assign w42479 = w42503 ^ w42474;
	assign w50871 = w45152 ^ w42479;
	assign w10467 = w50871 ^ w50876;
	assign w10309 = ~w10467;
	assign w10306 = w10309 ^ w10464;
	assign w50781 = w10306 ^ w10307;
	assign w46168 = w50781 ^ w699;
	assign w2982 = w46170 ^ w46168;
	assign w2980 = w46168 ^ w46165;
	assign w10332 = w10467 ^ w10454;
	assign w50773 = w10520 ^ w10467;
	assign w46176 = w50773 ^ w691;
	assign w42284 = w46178 ^ w46176;
	assign w42282 = w46176 ^ w46173;
	assign w10351 = w45838 ^ w50871;
	assign w50758 = w10350 ^ w10351;
	assign w46191 = w50758 ^ w676;
	assign w42453 = w42496 ^ w42497;
	assign w42554 = w42479 ^ w42453;
	assign w45874 = ~w42556;
	assign w10194 = w40545 ^ w45874;
	assign w10527 = w10193 ^ w10194;
	assign w50754 = w10527 ^ w10472;
	assign w10479 = w45874 ^ w45840;
	assign w10318 = w10479 ^ w10438;
	assign w50777 = w45878 ^ w10318;
	assign w10340 = w10479 ^ w10472;
	assign w10328 = w10479 ^ w10446;
	assign w50769 = w45807 ^ w10328;
	assign w46172 = w50777 ^ w695;
	assign w46180 = w50769 ^ w687;
	assign w50761 = w45874 ^ w10342;
	assign w46188 = w50761 ^ w679;
	assign w46195 = w50754 ^ w672;
	assign w2623 = w46195 ^ w46193;
	assign w45879 = ~w42553;
	assign w10349 = w45812 ^ w45879;
	assign w50759 = w10348 ^ w10349;
	assign w46190 = w50759 ^ w677;
	assign w2626 = w46192 ^ w46190;
	assign w2630 = w46196 ^ w46190;
	assign w2585 = w2626 ^ w46191;
	assign w2709 = w46196 ^ w2585;
	assign w2695 = w46196 & w2709;
	assign w2710 = w46191 ^ w2630;
	assign w2706 = w46195 ^ w2710;
	assign w2693 = w2710 & w2706;
	assign w10463 = w45879 ^ w45838;
	assign w10324 = w10463 ^ w45812;
	assign w10322 = ~w10324;
	assign w50774 = w10322 ^ w10323;
	assign w46175 = w50774 ^ w692;
	assign w42194 = w46175 ^ w46173;
	assign w42269 = w42194 ^ w42284;
	assign w42260 = w42284 & w42269;
	assign w50766 = w45879 ^ w10332;
	assign w46183 = w50766 ^ w684;
	assign w10305 = w10463 ^ w10459;
	assign w50782 = w45883 ^ w10305;
	assign w46167 = w50782 ^ w700;
	assign w2892 = w46167 ^ w46165;
	assign w2967 = w2892 ^ w2982;
	assign w2958 = w2982 & w2967;
	assign w45880 = ~w42554;
	assign w50783 = w45880 ^ w10304;
	assign w46166 = w50783 ^ w701;
	assign w10330 = w50872 ^ w45880;
	assign w2894 = w46168 ^ w46166;
	assign w2853 = w2894 ^ w46167;
	assign w2977 = w46172 ^ w2853;
	assign w2898 = w46172 ^ w46166;
	assign w2975 = w2892 ^ w2898;
	assign w10457 = w45880 ^ w45813;
	assign w10320 = w10457 ^ w45883;
	assign w50775 = w10320 ^ w10321;
	assign w46174 = w50775 ^ w693;
	assign w42196 = w46176 ^ w46174;
	assign w42155 = w42196 ^ w46175;
	assign w42279 = w46180 ^ w42155;
	assign w42200 = w46180 ^ w46174;
	assign w42280 = w46175 ^ w42200;
	assign w50768 = w10329 ^ w10330;
	assign w46181 = w50768 ^ w686;
	assign w2758 = w46183 ^ w46181;
	assign w42156 = w42196 ^ w42194;
	assign w2963 = w46172 & w2977;
	assign w2854 = w2894 ^ w2892;
	assign w10347 = w10457 ^ w10438;
	assign w50760 = w50877 ^ w10347;
	assign w46189 = w50760 ^ w678;
	assign w2712 = w46192 ^ w46189;
	assign w2713 = w46189 ^ w46195;
	assign w2704 = w2623 ^ w2712;
	assign w2703 = w46196 ^ w2704;
	assign w2624 = w46191 ^ w46189;
	assign w2707 = w2624 ^ w2630;
	assign w2586 = w2626 ^ w2624;
	assign w2702 = w2623 ^ w2586;
	assign w42265 = w46180 & w42279;
	assign w2978 = w46167 ^ w2898;
	assign w45881 = ~w42555;
	assign w10478 = w45881 ^ w50873;
	assign w10353 = w50874 ^ w45881;
	assign w50755 = w10352 ^ w10353;
	assign w46194 = w50755 ^ w673;
	assign w2640 = w46195 ^ w46194;
	assign w2708 = w2712 ^ w2640;
	assign w2697 = w2704 & w2708;
	assign w2629 = w2697 ^ w2626;
	assign w2711 = w46189 ^ w46194;
	assign w2689 = w2711 & w2702;
	assign w43645 = w2689 ^ w2695;
	assign w2639 = w43645 ^ w2624;
	assign w10338 = w10478 ^ w10469;
	assign w10316 = w10478 ^ w10476;
	assign w50778 = w10316 ^ w10317;
	assign w46171 = w50778 ^ w696;
	assign w2974 = w46171 ^ w2978;
	assign w2891 = w46171 ^ w46169;
	assign w2981 = w46165 ^ w46171;
	assign w2961 = w2978 & w2974;
	assign w2893 = w46170 ^ w2891;
	assign w2966 = w46167 ^ w2893;
	assign w2969 = w46166 ^ w2893;
	assign w2968 = w2898 ^ w2893;
	assign w2960 = w2975 & w2968;
	assign w2962 = w2981 & w2966;
	assign w2896 = w2962 ^ w2892;
	assign w2970 = w2891 ^ w2854;
	assign w2957 = w2979 & w2970;
	assign w50763 = w50869 ^ w10338;
	assign w46186 = w50763 ^ w681;
	assign w2845 = w46181 ^ w46186;
	assign w2959 = w2980 & w2969;
	assign w2867 = w2958 ^ w2959;
	assign w50770 = w10522 ^ w10478;
	assign w46179 = w50770 ^ w688;
	assign w42193 = w46179 ^ w46177;
	assign w42210 = w46179 ^ w46178;
	assign w42274 = w42193 ^ w42282;
	assign w42195 = w46178 ^ w42193;
	assign w42270 = w42200 ^ w42195;
	assign w42276 = w46179 ^ w42280;
	assign w42263 = w42280 & w42276;
	assign w42271 = w46174 ^ w42195;
	assign w42261 = w42282 & w42271;
	assign w42197 = w42261 ^ w42195;
	assign w42169 = w42260 ^ w42261;
	assign w42216 = w42169 ^ w42170;
	assign w42268 = w46175 ^ w42195;
	assign w42278 = w42282 ^ w42210;
	assign w42267 = w42274 & w42278;
	assign w42199 = w42267 ^ w42196;
	assign w42203 = w42199 ^ w42197;
	assign w42208 = w46173 ^ w42203;
	assign w2625 = w46194 ^ w2623;
	assign w2700 = w2630 ^ w2625;
	assign w2698 = w46191 ^ w2625;
	assign w2692 = w2707 & w2700;
	assign w2694 = w2713 & w2698;
	assign w2628 = w2694 ^ w2624;
	assign w2701 = w46190 ^ w2625;
	assign w2691 = w2712 & w2701;
	assign w2627 = w2691 ^ w2625;
	assign w2714 = w46194 ^ w46192;
	assign w2699 = w2624 ^ w2714;
	assign w2690 = w2714 & w2699;
	assign w2599 = w2690 ^ w2691;
	assign w42283 = w46173 ^ w46179;
	assign w42264 = w42283 & w42268;
	assign w42198 = w42264 ^ w42194;
	assign w42273 = w46180 ^ w42274;
	assign w42215 = w42216 ^ w42198;
	assign w42257 = w42263 ^ w42215;
	assign w2633 = w2629 ^ w2627;
	assign w2601 = w2633 ^ w43645;
	assign w2644 = w46191 ^ w2601;
	assign w2638 = w46189 ^ w2633;
	assign w2972 = w2891 ^ w2980;
	assign w2971 = w46172 ^ w2972;
	assign w43653 = w2957 ^ w2963;
	assign w2907 = w43653 ^ w2892;
	assign w2895 = w2959 ^ w2893;
	assign w2600 = w46193 ^ w46194;
	assign w2646 = w2599 ^ w2600;
	assign w2645 = w2646 ^ w2628;
	assign w2687 = w2693 ^ w2645;
	assign w43642 = w2689 ^ w2692;
	assign w2642 = w2690 ^ w43642;
	assign w2598 = w2693 ^ w2642;
	assign w2602 = w2628 ^ w43642;
	assign w2686 = w2602 ^ w2627;
	assign w2680 = w46195 ^ w2598;
	assign w2908 = w46171 ^ w46170;
	assign w2976 = w2980 ^ w2908;
	assign w2973 = w2908 ^ w2975;
	assign w2965 = w2972 & w2976;
	assign w2897 = w2965 ^ w2894;
	assign w2901 = w2897 ^ w2895;
	assign w2906 = w46165 ^ w2901;
	assign w2869 = w2901 ^ w43653;
	assign w2964 = w2973 & w2971;
	assign w43654 = w2957 ^ w2960;
	assign w2910 = w2958 ^ w43654;
	assign w2866 = w2961 ^ w2910;
	assign w2948 = w46171 ^ w2866;
	assign w42272 = w42193 ^ w42156;
	assign w42259 = w42281 & w42272;
	assign w45139 = w42259 ^ w42265;
	assign w42209 = w45139 ^ w42194;
	assign w42171 = w42203 ^ w45139;
	assign w42214 = w46175 ^ w42171;
	assign w2870 = w2896 ^ w43654;
	assign w2954 = w2870 ^ w2895;
	assign w10331 = w10463 ^ w10457;
	assign w50767 = w45884 ^ w10331;
	assign w46182 = w50767 ^ w685;
	assign w2764 = w46188 ^ w46182;
	assign w2841 = w2758 ^ w2764;
	assign w2844 = w46183 ^ w2764;
	assign w2705 = w2640 ^ w2707;
	assign w2696 = w2705 & w2703;
	assign w2647 = w2690 ^ w2696;
	assign w2685 = w2647 ^ w2639;
	assign w2688 = w2647 ^ w2638;
	assign w2684 = w2688 & w2687;
	assign w2683 = w2684 ^ w2686;
	assign w2682 = w2685 & w2683;
	assign w2593 = w2682 ^ w2694;
	assign w2589 = w2593 ^ w2629;
	assign w2592 = w46189 ^ w2589;
	assign w2588 = w46191 ^ w2589;
	assign w2681 = w2682 ^ w2644;
	assign w2651 = w2681 & w2707;
	assign w2679 = w2684 ^ w2644;
	assign w2678 = w2679 & w2680;
	assign w2596 = w2678 ^ w2695;
	assign w2591 = w2596 ^ w2692;
	assign w2676 = w2684 ^ w2678;
	assign w2675 = w2686 & w2676;
	assign w2673 = w2675 ^ w2683;
	assign w2672 = w2681 & w2673;
	assign w2595 = w2672 ^ w2696;
	assign w2637 = w2672 ^ w2647;
	assign w2671 = w2637 ^ w2639;
	assign w2652 = w2671 & w2706;
	assign w2661 = w2671 & w2710;
	assign w43644 = w2675 ^ w2693;
	assign w2634 = w46195 ^ w43644;
	assign w2587 = w2634 ^ w2595;
	assign w2666 = w2587 ^ w2588;
	assign w2658 = w2666 & w2699;
	assign w2597 = w2678 ^ w2642;
	assign w2674 = w2634 ^ w2597;
	assign w2664 = w2674 & w2703;
	assign w2619 = w2658 ^ w2661;
	assign w2616 = ~w2619;
	assign w2649 = w2666 & w2714;
	assign w2677 = w2678 ^ w2686;
	assign w2654 = w2677 & w2709;
	assign w2663 = w2677 & w46196;
	assign w2590 = w2682 ^ w2638;
	assign w2668 = w2637 ^ w2590;
	assign w2662 = w2668 & w2698;
	assign w43646 = w2661 ^ w2662;
	assign w2653 = w2668 & w2713;
	assign w2620 = w2662 ^ w2653;
	assign w2594 = w2624 ^ w2587;
	assign w2670 = w2591 ^ w2594;
	assign w2648 = w2670 & w2711;
	assign w2657 = w2670 & w2702;
	assign w2635 = w2653 ^ w2657;
	assign w2613 = ~w2635;
	assign w2612 = w2613 ^ w2651;
	assign w2667 = w43644 ^ w2645;
	assign w2656 = w2667 & w2708;
	assign w2665 = w2667 & w2704;
	assign w43647 = w2663 ^ w2665;
	assign w2608 = w2612 ^ w43647;
	assign w2643 = w2658 ^ w43646;
	assign w2609 = w2654 ^ w2643;
	assign w2606 = ~w2609;
	assign w2660 = w2681 & w2700;
	assign w2604 = w2660 ^ w2661;
	assign w2622 = w2660 ^ w2652;
	assign w2669 = w2591 ^ w2592;
	assign w2650 = w2669 & w2712;
	assign w43643 = w2649 ^ w2650;
	assign w2618 = w2622 ^ w43643;
	assign w2617 = w2613 ^ w2618;
	assign w2717 = w2616 ^ w2617;
	assign w2659 = w2669 & w2701;
	assign w2603 = w2659 ^ w2643;
	assign w2615 = w2658 ^ w2659;
	assign w2614 = w2659 ^ w2648;
	assign w2610 = ~w2614;
	assign w2621 = w43647 ^ w2618;
	assign w45974 = ~w2717;
	assign w50923 = w45974 ^ w832;
	assign w2611 = w2650 ^ w2608;
	assign w2715 = w2610 ^ w2611;
	assign w45978 = ~w2715;
	assign w50927 = w45978 ^ w836;
	assign w2655 = w2674 & w2705;
	assign w2631 = w2655 ^ w43643;
	assign w2632 = w2656 ^ w2631;
	assign w45980 = w2632 ^ w2603;
	assign w50929 = w45980 ^ w838;
	assign w2636 = w2664 ^ w2632;
	assign w2605 = w2663 ^ w2636;
	assign w45976 = w2604 ^ w2605;
	assign w2641 = w2665 ^ w2636;
	assign w50925 = w45976 ^ w834;
	assign w2716 = w2641 ^ w2615;
	assign w45979 = ~w2716;
	assign w50928 = w45979 ^ w837;
	assign w2607 = w2631 ^ w2608;
	assign w45975 = w2606 ^ w2607;
	assign w50924 = w45975 ^ w833;
	assign w2915 = w2958 ^ w2964;
	assign w2953 = w2915 ^ w2907;
	assign w2956 = w2915 ^ w2906;
	assign w2127 = w2141 & w46228;
	assign w43623 = w2127 ^ w2129;
	assign w2088 = w2084 ^ w43623;
	assign w2085 = w2114 ^ w2088;
	assign w2179 = w2086 ^ w2085;
	assign w46074 = ~w2179;
	assign w51023 = w46074 ^ w740;
	assign w2089 = w2065 ^ w2088;
	assign w46071 = w2090 ^ w2089;
	assign w51020 = w46071 ^ w737;
	assign w2075 = w43623 ^ w2078;
	assign w2182 = w2076 ^ w2075;
	assign w46069 = ~w2182;
	assign w51018 = w46069 ^ w735;
	assign w2718 = w2620 ^ w2621;
	assign w45973 = ~w2718;
	assign w50922 = w45973 ^ w831;
	assign w2120 = w2131 & w2172;
	assign w2064 = w2120 ^ w2065;
	assign w2059 = w2128 ^ w2064;
	assign w2054 = w2129 ^ w2059;
	assign w2180 = w2054 ^ w2081;
	assign w46076 = w2064 ^ w2093;
	assign w46073 = w43622 ^ w2054;
	assign w2091 = w2127 ^ w2059;
	assign w51022 = w46073 ^ w739;
	assign w46072 = w2092 ^ w2091;
	assign w51021 = w46072 ^ w738;
	assign w51025 = w46076 ^ w742;
	assign w46075 = ~w2180;
	assign w51024 = w46075 ^ w741;
	assign w45977 = w43646 ^ w2641;
	assign w50926 = w45977 ^ w835;
	assign w50614 = w45834 ^ w9635;
	assign w46262 = w50614 ^ w541;
	assign w39859 = w46262 ^ w39783;
	assign w39784 = w46264 ^ w46262;
	assign w39787 = w39855 ^ w39784;
	assign w39743 = w39784 ^ w46263;
	assign w39744 = w39784 ^ w39782;
	assign w39849 = w39870 & w39859;
	assign w39785 = w39849 ^ w39783;
	assign w39791 = w39787 ^ w39785;
	assign w39796 = w46261 ^ w39791;
	assign w39757 = w39848 ^ w39849;
	assign w39804 = w39757 ^ w39758;
	assign w39803 = w39804 ^ w39786;
	assign w42277 = w42194 ^ w42200;
	assign w42262 = w42277 & w42270;
	assign w45140 = w42259 ^ w42262;
	assign w42212 = w42260 ^ w45140;
	assign w42168 = w42263 ^ w42212;
	assign w42250 = w46179 ^ w42168;
	assign w42275 = w42210 ^ w42277;
	assign w42266 = w42275 & w42273;
	assign w42217 = w42260 ^ w42266;
	assign w42258 = w42217 ^ w42208;
	assign w42254 = w42258 & w42257;
	assign w42249 = w42254 ^ w42214;
	assign w42248 = w42249 & w42250;
	assign w42246 = w42254 ^ w42248;
	assign w42255 = w42217 ^ w42209;
	assign w42167 = w42248 ^ w42212;
	assign w42172 = w42198 ^ w45140;
	assign w42256 = w42172 ^ w42197;
	assign w42247 = w42248 ^ w42256;
	assign w42233 = w42247 & w46180;
	assign w42253 = w42254 ^ w42256;
	assign w42245 = w42256 & w42246;
	assign w45143 = w42245 ^ w42263;
	assign w42204 = w46179 ^ w45143;
	assign w42244 = w42204 ^ w42167;
	assign w42234 = w42244 & w42273;
	assign w42237 = w45143 ^ w42215;
	assign w42226 = w42237 & w42278;
	assign w42252 = w42255 & w42253;
	assign w42163 = w42252 ^ w42264;
	assign w42160 = w42252 ^ w42208;
	assign w42251 = w42252 ^ w42214;
	assign w42221 = w42251 & w42277;
	assign w42230 = w42251 & w42270;
	assign w42235 = w42237 & w42274;
	assign w45142 = w42233 ^ w42235;
	assign w42243 = w42245 ^ w42253;
	assign w42242 = w42251 & w42243;
	assign w42207 = w42242 ^ w42217;
	assign w42238 = w42207 ^ w42160;
	assign w42241 = w42207 ^ w42209;
	assign w42232 = w42238 & w42268;
	assign w42165 = w42242 ^ w42266;
	assign w42157 = w42204 ^ w42165;
	assign w42164 = w42194 ^ w42157;
	assign w42223 = w42238 & w42283;
	assign w42222 = w42241 & w42276;
	assign w42231 = w42241 & w42280;
	assign w45141 = w42231 ^ w42232;
	assign w42225 = w42244 & w42275;
	assign w42174 = w42230 ^ w42231;
	assign w42224 = w42247 & w42279;
	assign w42166 = w42248 ^ w42265;
	assign w42161 = w42166 ^ w42262;
	assign w42240 = w42161 ^ w42164;
	assign w42227 = w42240 & w42272;
	assign w42218 = w42240 & w42281;
	assign w42159 = w42163 ^ w42199;
	assign w42158 = w46175 ^ w42159;
	assign w42236 = w42157 ^ w42158;
	assign w42228 = w42236 & w42269;
	assign w42219 = w42236 & w42284;
	assign w42162 = w46173 ^ w42159;
	assign w42239 = w42161 ^ w42162;
	assign w42220 = w42239 & w42282;
	assign w43616 = w42219 ^ w42220;
	assign w42201 = w42225 ^ w43616;
	assign w42229 = w42239 & w42271;
	assign w42184 = w42229 ^ w42218;
	assign w42180 = ~w42184;
	assign w42185 = w42228 ^ w42229;
	assign w42213 = w42228 ^ w45141;
	assign w42173 = w42229 ^ w42213;
	assign w42179 = w42224 ^ w42213;
	assign w42176 = ~w42179;
	assign w42202 = w42226 ^ w42201;
	assign w46060 = w42202 ^ w42173;
	assign w51009 = w46060 ^ w790;
	assign w42206 = w42234 ^ w42202;
	assign w42211 = w42235 ^ w42206;
	assign w46057 = w45141 ^ w42211;
	assign w51006 = w46057 ^ w787;
	assign w42189 = w42228 ^ w42231;
	assign w42186 = ~w42189;
	assign w42175 = w42233 ^ w42206;
	assign w46056 = w42174 ^ w42175;
	assign w51005 = w46056 ^ w786;
	assign w42286 = w42211 ^ w42185;
	assign w46059 = ~w42286;
	assign w51008 = w46059 ^ w789;
	assign w42205 = w42223 ^ w42227;
	assign w42183 = ~w42205;
	assign w42182 = w42183 ^ w42221;
	assign w42178 = w42182 ^ w45142;
	assign w42181 = w42220 ^ w42178;
	assign w42285 = w42180 ^ w42181;
	assign w42177 = w42201 ^ w42178;
	assign w46055 = w42176 ^ w42177;
	assign w46058 = ~w42285;
	assign w51007 = w46058 ^ w788;
	assign w51004 = w46055 ^ w785;
	assign w42192 = w42230 ^ w42222;
	assign w42188 = w42192 ^ w43616;
	assign w42187 = w42183 ^ w42188;
	assign w42191 = w45142 ^ w42188;
	assign w42287 = w42186 ^ w42187;
	assign w46054 = ~w42287;
	assign w51003 = w46054 ^ w784;
	assign w10380 = w10504 ^ w10482;
	assign w10379 = w10380 ^ w10381;
	assign w50738 = ~w10379;
	assign w46211 = w50738 ^ w720;
	assign w2355 = w46211 ^ w46209;
	assign w2357 = w46210 ^ w2355;
	assign w2430 = w46207 ^ w2357;
	assign w2432 = w2362 ^ w2357;
	assign w2433 = w46206 ^ w2357;
	assign w2372 = w46211 ^ w46210;
	assign w2438 = w46211 ^ w2442;
	assign w2425 = w2442 & w2438;
	assign w9648 = w9890 ^ w9824;
	assign w50608 = w45836 ^ w9648;
	assign w46268 = w50608 ^ w535;
	assign w39867 = w46268 ^ w39743;
	assign w39788 = w46268 ^ w46262;
	assign w39865 = w39782 ^ w39788;
	assign w39858 = w39788 ^ w39783;
	assign w39868 = w46263 ^ w39788;
	assign w39864 = w46267 ^ w39868;
	assign w39851 = w39868 & w39864;
	assign w39853 = w46268 & w39867;
	assign w39845 = w39851 ^ w39803;
	assign w39863 = w39798 ^ w39865;
	assign w39861 = w46268 ^ w39862;
	assign w39854 = w39863 & w39861;
	assign w39805 = w39848 ^ w39854;
	assign w39846 = w39805 ^ w39796;
	assign w39842 = w39846 & w39845;
	assign w39850 = w39865 & w39858;
	assign w41265 = w41261 ^ w41259;
	assign w41270 = w46269 ^ w41265;
	assign w39860 = w39781 ^ w39744;
	assign w39847 = w39869 & w39860;
	assign w45041 = w39847 ^ w39853;
	assign w39797 = w45041 ^ w39782;
	assign w39843 = w39805 ^ w39797;
	assign w39759 = w39791 ^ w45041;
	assign w39802 = w46263 ^ w39759;
	assign w39837 = w39842 ^ w39802;
	assign w45038 = w39847 ^ w39850;
	assign w39800 = w39848 ^ w45038;
	assign w39756 = w39851 ^ w39800;
	assign w39838 = w46267 ^ w39756;
	assign w39836 = w39837 & w39838;
	assign w39834 = w39842 ^ w39836;
	assign w39755 = w39836 ^ w39800;
	assign w39754 = w39836 ^ w39853;
	assign w39749 = w39754 ^ w39850;
	assign w39760 = w39786 ^ w45038;
	assign w39844 = w39760 ^ w39785;
	assign w39833 = w39844 & w39834;
	assign w39835 = w39836 ^ w39844;
	assign w39821 = w39835 & w46268;
	assign w45040 = w39833 ^ w39851;
	assign w39825 = w45040 ^ w39803;
	assign w39823 = w39825 & w39862;
	assign w45043 = w39821 ^ w39823;
	assign w39841 = w39842 ^ w39844;
	assign w39792 = w46267 ^ w45040;
	assign w39832 = w39792 ^ w39755;
	assign w39814 = w39825 & w39866;
	assign w39840 = w39843 & w39841;
	assign w39748 = w39840 ^ w39796;
	assign w39839 = w39840 ^ w39802;
	assign w39818 = w39839 & w39858;
	assign w39822 = w39832 & w39861;
	assign w39751 = w39840 ^ w39852;
	assign w39747 = w39751 ^ w39787;
	assign w39750 = w46261 ^ w39747;
	assign w39831 = w39833 ^ w39841;
	assign w39830 = w39839 & w39831;
	assign w39753 = w39830 ^ w39854;
	assign w39745 = w39792 ^ w39753;
	assign w39752 = w39782 ^ w39745;
	assign w39828 = w39749 ^ w39752;
	assign w39806 = w39828 & w39869;
	assign w39815 = w39828 & w39860;
	assign w39795 = w39830 ^ w39805;
	assign w39829 = w39795 ^ w39797;
	assign w39826 = w39795 ^ w39748;
	assign w39811 = w39826 & w39871;
	assign w39819 = w39829 & w39868;
	assign w39762 = w39818 ^ w39819;
	assign w39793 = w39811 ^ w39815;
	assign w39810 = w39829 & w39864;
	assign w39780 = w39818 ^ w39810;
	assign w39820 = w39826 & w39856;
	assign w39778 = w39820 ^ w39811;
	assign w39812 = w39835 & w39867;
	assign w45042 = w39819 ^ w39820;
	assign w39771 = ~w39793;
	assign w39827 = w39749 ^ w39750;
	assign w39808 = w39827 & w39870;
	assign w39817 = w39827 & w39859;
	assign w39772 = w39817 ^ w39806;
	assign w39768 = ~w39772;
	assign w39813 = w39832 & w39863;
	assign w39746 = w46263 ^ w39747;
	assign w39824 = w39745 ^ w39746;
	assign w39807 = w39824 & w39872;
	assign w45039 = w39807 ^ w39808;
	assign w39789 = w39813 ^ w45039;
	assign w39776 = w39780 ^ w45039;
	assign w39779 = w45043 ^ w39776;
	assign w39775 = w39771 ^ w39776;
	assign w39876 = w39778 ^ w39779;
	assign w39790 = w39814 ^ w39789;
	assign w39794 = w39822 ^ w39790;
	assign w39799 = w39823 ^ w39794;
	assign w39763 = w39821 ^ w39794;
	assign w50902 = w39762 ^ w39763;
	assign w50903 = w45042 ^ w39799;
	assign w10226 = w10225 ^ w50903;
	assign w10477 = w50898 ^ w50902;
	assign w10250 = w10252 ^ w10477;
	assign w10280 = w10271 ^ w10477;
	assign w50796 = w10280 ^ w10281;
	assign w46153 = w50796 ^ w650;
	assign w10514 = w10226 ^ w10227;
	assign w50805 = w10514 ^ w10480;
	assign w46144 = w50805 ^ w659;
	assign w39816 = w39824 & w39857;
	assign w39773 = w39816 ^ w39817;
	assign w39874 = w39799 ^ w39773;
	assign w39801 = w39816 ^ w45042;
	assign w39767 = w39812 ^ w39801;
	assign w39764 = ~w39767;
	assign w10222 = w10225 ^ w50902;
	assign w10515 = w10222 ^ w10223;
	assign w50804 = w10515 ^ w10488;
	assign w46145 = w50804 ^ w658;
	assign w10468 = w50899 ^ w50903;
	assign w10278 = w10255 ^ w10468;
	assign w50797 = w10278 ^ w10279;
	assign w46152 = w50797 ^ w651;
	assign w10249 = w10473 ^ w10468;
	assign w50814 = w45860 ^ w10249;
	assign w46135 = w50814 ^ w668;
	assign w45822 = ~w39874;
	assign w10266 = w10466 ^ w45822;
	assign w10264 = ~w10266;
	assign w50807 = w10264 ^ w10265;
	assign w46142 = w50807 ^ w661;
	assign w40320 = w46144 ^ w46142;
	assign w10451 = w45861 ^ w45822;
	assign w10247 = w10451 ^ w10440;
	assign w50816 = w50900 ^ w10247;
	assign w46133 = w50816 ^ w670;
	assign w39648 = w46135 ^ w46133;
	assign w10276 = w10473 ^ w10451;
	assign w50799 = w45853 ^ w10276;
	assign w46150 = w50799 ^ w653;
	assign w40990 = w46152 ^ w46150;
	assign w45824 = ~w39876;
	assign w50801 = w45824 ^ w10272;
	assign w46148 = w50801 ^ w655;
	assign w40324 = w46148 ^ w46142;
	assign w10499 = w45855 ^ w45824;
	assign w10286 = w10499 ^ w10440;
	assign w50793 = w45847 ^ w10286;
	assign w46156 = w50793 ^ w647;
	assign w39761 = w39817 ^ w39801;
	assign w50904 = w39790 ^ w39761;
	assign w10437 = w50900 ^ w50904;
	assign w10275 = w10466 ^ w10437;
	assign w50800 = w50889 ^ w10275;
	assign w10261 = w10503 ^ w10437;
	assign w46149 = w50800 ^ w654;
	assign w41076 = w46152 ^ w46149;
	assign w10287 = w10437 ^ w45822;
	assign w50792 = w10287 ^ w10288;
	assign w46157 = w50792 ^ w646;
	assign w10262 = w45894 ^ w50904;
	assign w50808 = w10262 ^ w10263;
	assign w46141 = w50808 ^ w662;
	assign w40406 = w46144 ^ w46141;
	assign w10445 = w50889 ^ w50904;
	assign w10218 = w10445 ^ w50902;
	assign w10517 = w10218 ^ w10219;
	assign w50789 = w10517 ^ w10468;
	assign w46160 = w50789 ^ w643;
	assign w10301 = w10499 ^ w10445;
	assign w50785 = w45843 ^ w10301;
	assign w42148 = w46160 ^ w46157;
	assign w46164 = w50785 ^ w639;
	assign w10214 = ~w10445;
	assign w50809 = w45855 ^ w10261;
	assign w46140 = w50809 ^ w663;
	assign w10212 = w10214 ^ w45824;
	assign w10519 = w10212 ^ w10213;
	assign w40994 = w46156 ^ w46150;
	assign w10260 = w10502 ^ w10499;
	assign w10258 = ~w10260;
	assign w39777 = w39816 ^ w39819;
	assign w39774 = ~w39777;
	assign w39875 = w39774 ^ w39775;
	assign w45823 = ~w39875;
	assign w10220 = w10444 ^ w45823;
	assign w10491 = w45854 ^ w45823;
	assign w10256 = w10495 ^ w10491;
	assign w50786 = w10519 ^ w10491;
	assign w50811 = w50897 ^ w10256;
	assign w46138 = w50811 ^ w665;
	assign w39735 = w46133 ^ w46138;
	assign w46163 = w50786 ^ w640;
	assign w42149 = w46157 ^ w46163;
	assign w10516 = w10220 ^ w10221;
	assign w50802 = w10516 ^ w10502;
	assign w46147 = w50802 ^ w656;
	assign w40317 = w46147 ^ w46145;
	assign w40398 = w40317 ^ w40406;
	assign w40397 = w46148 ^ w40398;
	assign w40407 = w46141 ^ w46147;
	assign w10284 = w10503 ^ w10491;
	assign w10283 = w10284 ^ w10285;
	assign w50794 = ~w10283;
	assign w46155 = w50794 ^ w648;
	assign w40987 = w46155 ^ w46153;
	assign w41068 = w40987 ^ w41076;
	assign w41067 = w46156 ^ w41068;
	assign w41077 = w46149 ^ w46155;
	assign w45957 = ~w10439;
	assign w10334 = w45957 ^ w50871;
	assign w50765 = w10333 ^ w10334;
	assign w46184 = w50765 ^ w683;
	assign w2846 = w46184 ^ w46181;
	assign w2760 = w46184 ^ w46182;
	assign w10341 = w45957 ^ w45881;
	assign w10339 = w10340 ^ w10341;
	assign w10337 = w45957 ^ w50870;
	assign w50764 = w10336 ^ w10337;
	assign w46185 = w50764 ^ w682;
	assign w2734 = w46185 ^ w46186;
	assign w2719 = w2760 ^ w46183;
	assign w2843 = w46188 ^ w2719;
	assign w2829 = w46188 & w2843;
	assign w2848 = w46186 ^ w46184;
	assign w2833 = w2758 ^ w2848;
	assign w2824 = w2848 & w2833;
	assign w50762 = ~w10339;
	assign w46187 = w50762 ^ w680;
	assign w2847 = w46181 ^ w46187;
	assign w2757 = w46187 ^ w46185;
	assign w2759 = w46186 ^ w2757;
	assign w2835 = w46182 ^ w2759;
	assign w2832 = w46183 ^ w2759;
	assign w2828 = w2847 & w2832;
	assign w2762 = w2828 ^ w2758;
	assign w2834 = w2764 ^ w2759;
	assign w2825 = w2846 & w2835;
	assign w2733 = w2824 ^ w2825;
	assign w2761 = w2825 ^ w2759;
	assign w2780 = w2733 ^ w2734;
	assign w2779 = w2780 ^ w2762;
	assign w2774 = w46187 ^ w46186;
	assign w2840 = w46187 ^ w2844;
	assign w2827 = w2844 & w2840;
	assign w2821 = w2827 ^ w2779;
	assign w2842 = w2846 ^ w2774;
	assign w2838 = w2757 ^ w2846;
	assign w2831 = w2838 & w2842;
	assign w2763 = w2831 ^ w2760;
	assign w2837 = w46188 ^ w2838;
	assign w2767 = w2763 ^ w2761;
	assign w2839 = w2774 ^ w2841;
	assign w2830 = w2839 & w2837;
	assign w2781 = w2824 ^ w2830;
	assign w2772 = w46181 ^ w2767;
	assign w2822 = w2781 ^ w2772;
	assign w2818 = w2822 & w2821;
	assign w2826 = w2841 & w2834;
	assign w2720 = w2760 ^ w2758;
	assign w2836 = w2757 ^ w2720;
	assign w2823 = w2845 & w2836;
	assign w43648 = w2823 ^ w2829;
	assign w2773 = w43648 ^ w2758;
	assign w2819 = w2781 ^ w2773;
	assign w2735 = w2767 ^ w43648;
	assign w2778 = w46183 ^ w2735;
	assign w2813 = w2818 ^ w2778;
	assign w45958 = ~w10437;
	assign w10251 = w45958 ^ w50899;
	assign w50813 = w10250 ^ w10251;
	assign w46136 = w50813 ^ w667;
	assign w39736 = w46136 ^ w46133;
	assign w10259 = w45958 ^ w45854;
	assign w50810 = w10258 ^ w10259;
	assign w46139 = w50810 ^ w664;
	assign w39664 = w46139 ^ w46138;
	assign w39732 = w39736 ^ w39664;
	assign w39737 = w46133 ^ w46139;
	assign w39738 = w46138 ^ w46136;
	assign w39723 = w39648 ^ w39738;
	assign w39714 = w39738 & w39723;
	assign w10254 = w45958 ^ w50898;
	assign w50600 = w45816 ^ w9659;
	assign w46276 = w50600 ^ w527;
	assign w41335 = w46276 ^ w41336;
	assign w41262 = w46276 ^ w46270;
	assign w41339 = w41256 ^ w41262;
	assign w41332 = w41262 ^ w41257;
	assign w41324 = w41339 & w41332;
	assign w41337 = w41272 ^ w41339;
	assign w41328 = w41337 & w41335;
	assign w45100 = w41321 ^ w41324;
	assign w41274 = w41322 ^ w45100;
	assign w41234 = w41260 ^ w45100;
	assign w41318 = w41234 ^ w41259;
	assign w41341 = w46276 ^ w41217;
	assign w41327 = w46276 & w41341;
	assign w41279 = w41322 ^ w41328;
	assign w41320 = w41279 ^ w41270;
	assign w45103 = w41321 ^ w41327;
	assign w41271 = w45103 ^ w41256;
	assign w41317 = w41279 ^ w41271;
	assign w41233 = w41265 ^ w45103;
	assign w41276 = w46271 ^ w41233;
	assign w41342 = w46271 ^ w41262;
	assign w41338 = w46275 ^ w41342;
	assign w41325 = w41342 & w41338;
	assign w41230 = w41325 ^ w41274;
	assign w41312 = w46275 ^ w41230;
	assign w41319 = w41325 ^ w41277;
	assign w41316 = w41320 & w41319;
	assign w41311 = w41316 ^ w41276;
	assign w41310 = w41311 & w41312;
	assign w41229 = w41310 ^ w41274;
	assign w41228 = w41310 ^ w41327;
	assign w41223 = w41228 ^ w41324;
	assign w41315 = w41316 ^ w41318;
	assign w41314 = w41317 & w41315;
	assign w41225 = w41314 ^ w41326;
	assign w41222 = w41314 ^ w41270;
	assign w41313 = w41314 ^ w41276;
	assign w41292 = w41313 & w41332;
	assign w41309 = w41310 ^ w41318;
	assign w41286 = w41309 & w41341;
	assign w41295 = w41309 & w46276;
	assign w41283 = w41313 & w41339;
	assign w41308 = w41316 ^ w41310;
	assign w41307 = w41318 & w41308;
	assign w45102 = w41307 ^ w41325;
	assign w41299 = w45102 ^ w41277;
	assign w41266 = w46275 ^ w45102;
	assign w41306 = w41266 ^ w41229;
	assign w41287 = w41306 & w41337;
	assign w41305 = w41307 ^ w41315;
	assign w41304 = w41313 & w41305;
	assign w41269 = w41304 ^ w41279;
	assign w41227 = w41304 ^ w41328;
	assign w41303 = w41269 ^ w41271;
	assign w41284 = w41303 & w41338;
	assign w41254 = w41292 ^ w41284;
	assign w41293 = w41303 & w41342;
	assign w41219 = w41266 ^ w41227;
	assign w41226 = w41256 ^ w41219;
	assign w41302 = w41223 ^ w41226;
	assign w41280 = w41302 & w41343;
	assign w41289 = w41302 & w41334;
	assign w41300 = w41269 ^ w41222;
	assign w41285 = w41300 & w41345;
	assign w41267 = w41285 ^ w41289;
	assign w41245 = ~w41267;
	assign w41244 = w41245 ^ w41283;
	assign w41288 = w41299 & w41340;
	assign w41297 = w41299 & w41336;
	assign w45105 = w41295 ^ w41297;
	assign w41240 = w41244 ^ w45105;
	assign w41296 = w41306 & w41335;
	assign w41294 = w41300 & w41330;
	assign w45104 = w41293 ^ w41294;
	assign w41252 = w41294 ^ w41285;
	assign w41236 = w41292 ^ w41293;
	assign w41221 = w41225 ^ w41261;
	assign w41224 = w46269 ^ w41221;
	assign w41220 = w46271 ^ w41221;
	assign w41298 = w41219 ^ w41220;
	assign w41290 = w41298 & w41331;
	assign w41275 = w41290 ^ w45104;
	assign w41241 = w41286 ^ w41275;
	assign w41238 = ~w41241;
	assign w41281 = w41298 & w41346;
	assign w41251 = w41290 ^ w41293;
	assign w41248 = ~w41251;
	assign w41301 = w41223 ^ w41224;
	assign w41291 = w41301 & w41333;
	assign w41235 = w41291 ^ w41275;
	assign w41247 = w41290 ^ w41291;
	assign w41282 = w41301 & w41344;
	assign w45101 = w41281 ^ w41282;
	assign w41263 = w41287 ^ w45101;
	assign w41239 = w41263 ^ w41240;
	assign w41264 = w41288 ^ w41263;
	assign w41268 = w41296 ^ w41264;
	assign w41273 = w41297 ^ w41268;
	assign w50916 = w45104 ^ w41273;
	assign w10452 = w50916 ^ w50920;
	assign w10432 = w10461 ^ w10452;
	assign w50821 = w10432 ^ w10433;
	assign w46128 = w50821 ^ w611;
	assign w10404 = w10470 ^ w50916;
	assign w50838 = w10404 ^ w10405;
	assign w50829 = w10508 ^ w10452;
	assign w46120 = w50829 ^ w619;
	assign w41237 = w41295 ^ w41268;
	assign w50915 = w41236 ^ w41237;
	assign w10243 = w50916 ^ w50915;
	assign w10419 = w45959 ^ w50915;
	assign w50828 = w10418 ^ w10419;
	assign w46121 = w50828 ^ w618;
	assign w41243 = w41282 ^ w41240;
	assign w46111 = w50838 ^ w628;
	assign w50917 = w41264 ^ w41235;
	assign w10435 = w50917 ^ w50921;
	assign w10411 = w10500 ^ w10435;
	assign w50832 = w50909 ^ w10411;
	assign w10400 = w10498 ^ w10435;
	assign w46117 = w50832 ^ w622;
	assign w3248 = w46120 ^ w46117;
	assign w41348 = w41273 ^ w41247;
	assign w10455 = w50911 ^ w50915;
	assign w50820 = w10523 ^ w10455;
	assign w10406 = w10501 ^ w10455;
	assign w46129 = w50820 ^ w610;
	assign w50914 = w41238 ^ w41239;
	assign w10453 = w50914 ^ w50918;
	assign w10244 = w10453 ^ w45858;
	assign w50819 = w10244 ^ w10245;
	assign w46130 = w50819 ^ w609;
	assign w3116 = w46130 ^ w46128;
	assign w10421 = w10490 ^ w10453;
	assign w50827 = w50905 ^ w10421;
	assign w46122 = w50827 ^ w617;
	assign w3250 = w46122 ^ w46120;
	assign w3247 = w46117 ^ w46122;
	assign w3002 = w46129 ^ w46130;
	assign w3136 = w46121 ^ w46122;
	assign w10450 = w50913 ^ w50917;
	assign w10410 = w10498 ^ w10450;
	assign w50833 = w45803 ^ w10410;
	assign w10407 = w10450 ^ w50920;
	assign w10189 = w10450 ^ w50914;
	assign w10529 = w10189 ^ w10190;
	assign w50836 = w10529 ^ w10461;
	assign w10394 = w10455 ^ w10453;
	assign w41246 = w41291 ^ w41280;
	assign w41242 = ~w41246;
	assign w41347 = w41242 ^ w41243;
	assign w46116 = w50833 ^ w623;
	assign w50837 = w10406 ^ w10407;
	assign w46112 = w50837 ^ w627;
	assign w41250 = w41254 ^ w45101;
	assign w41249 = w41245 ^ w41250;
	assign w41349 = w41248 ^ w41249;
	assign w46113 = w50836 ^ w626;
	assign w10187 = w10450 ^ w45802;
	assign w10242 = w10435 ^ w50919;
	assign w10507 = w10242 ^ w10243;
	assign w50845 = w10507 ^ w10501;
	assign w46104 = w50845 ^ w635;
	assign w45850 = ~w41349;
	assign w10465 = w45850 ^ w45802;
	assign w10396 = w10475 ^ w10465;
	assign w50843 = w50914 ^ w10396;
	assign w10409 = w45850 ^ w45209;
	assign w46106 = w50843 ^ w633;
	assign w3518 = w46106 ^ w46104;
	assign w10423 = w10498 ^ w10465;
	assign w50818 = w10524 ^ w10465;
	assign w46131 = w50818 ^ w608;
	assign w3025 = w46131 ^ w46129;
	assign w3042 = w46131 ^ w46130;
	assign w3027 = w46130 ^ w3025;
	assign w45856 = ~w41347;
	assign w50830 = w45856 ^ w10417;
	assign w46119 = w50830 ^ w620;
	assign w3160 = w46119 ^ w46117;
	assign w3235 = w3160 ^ w3250;
	assign w10460 = w45212 ^ w45856;
	assign w10392 = w10460 ^ w10452;
	assign w50846 = w45865 ^ w10392;
	assign w46103 = w50846 ^ w636;
	assign w3226 = w3250 & w3235;
	assign w10403 = w10500 ^ w10460;
	assign w10431 = ~w10460;
	assign w10429 = w10431 ^ w45808;
	assign w50822 = w10429 ^ w10430;
	assign w46127 = w50822 ^ w612;
	assign w3100 = w46127 ^ w3027;
	assign w45857 = ~w41348;
	assign w10458 = w45857 ^ w45809;
	assign w10413 = w10458 ^ w45212;
	assign w10412 = w10413 ^ w10414;
	assign w10391 = w45857 ^ w45856;
	assign w10389 = w10458 ^ w10436;
	assign w50848 = w50917 ^ w10389;
	assign w46101 = w50848 ^ w638;
	assign w3516 = w46104 ^ w46101;
	assign w3515 = w46101 ^ w46106;
	assign w10428 = w10470 ^ w10458;
	assign w50823 = w45208 ^ w10428;
	assign w46126 = w50823 ^ w613;
	assign w3028 = w46128 ^ w46126;
	assign w50831 = ~w10412;
	assign w46118 = w50831 ^ w621;
	assign w3103 = w46126 ^ w3027;
	assign w3162 = w46120 ^ w46118;
	assign w50847 = w10390 ^ w10391;
	assign w46102 = w50847 ^ w637;
	assign w3428 = w46103 ^ w46101;
	assign w3503 = w3428 ^ w3518;
	assign w3494 = w3518 & w3503;
	assign w3430 = w46104 ^ w46102;
	assign w3390 = w3430 ^ w3428;
	assign w3389 = w3430 ^ w46103;
	assign w2987 = w3028 ^ w46127;
	assign w10402 = w45857 ^ w45208;
	assign w50840 = w10401 ^ w10402;
	assign w46109 = w50840 ^ w630;
	assign w3382 = w46112 ^ w46109;
	assign w3121 = w3162 ^ w46119;
	assign w3122 = w3162 ^ w3160;
	assign w3294 = w46111 ^ w46109;
	assign w41253 = w45105 ^ w41250;
	assign w41350 = w41252 ^ w41253;
	assign w45851 = ~w41350;
	assign w50841 = w45851 ^ w10400;
	assign w46108 = w50841 ^ w631;
	assign w3434 = w46108 ^ w46102;
	assign w3511 = w3428 ^ w3434;
	assign w3513 = w46108 ^ w3389;
	assign w3499 = w46108 & w3513;
	assign w3514 = w46103 ^ w3434;
	assign w10485 = w45851 ^ w45803;
	assign w10425 = w10485 ^ w10436;
	assign w10397 = w10399 ^ w10485;
	assign w10246 = w10485 ^ w10447;
	assign w50817 = w45210 ^ w10246;
	assign w46132 = w50817 ^ w607;
	assign w3111 = w46132 ^ w2987;
	assign w3097 = w46132 & w3111;
	assign w3032 = w46132 ^ w46126;
	assign w3102 = w3032 ^ w3027;
	assign w3112 = w46127 ^ w3032;
	assign w3108 = w46131 ^ w3112;
	assign w3095 = w3112 & w3108;
	assign w50825 = w45859 ^ w10425;
	assign w46124 = w50825 ^ w615;
	assign w3245 = w46124 ^ w3121;
	assign w3231 = w46124 & w3245;
	assign w3166 = w46124 ^ w46118;
	assign w3246 = w46119 ^ w3166;
	assign w3243 = w3160 ^ w3166;
	assign w10422 = w10423 ^ w10424;
	assign w50826 = ~w10422;
	assign w46123 = w50826 ^ w616;
	assign w3249 = w46117 ^ w46123;
	assign w3242 = w46123 ^ w3246;
	assign w3229 = w3246 & w3242;
	assign w3159 = w46123 ^ w46121;
	assign w3238 = w3159 ^ w3122;
	assign w3240 = w3159 ^ w3248;
	assign w3176 = w46123 ^ w46122;
	assign w3241 = w3176 ^ w3243;
	assign w3244 = w3248 ^ w3176;
	assign w3233 = w3240 & w3244;
	assign w3165 = w3233 ^ w3162;
	assign w3161 = w46122 ^ w3159;
	assign w3237 = w46118 ^ w3161;
	assign w3227 = w3248 & w3237;
	assign w3135 = w3226 ^ w3227;
	assign w3182 = w3135 ^ w3136;
	assign w3163 = w3227 ^ w3161;
	assign w3169 = w3165 ^ w3163;
	assign w3174 = w46117 ^ w3169;
	assign w3234 = w46119 ^ w3161;
	assign w3230 = w3249 & w3234;
	assign w3164 = w3230 ^ w3160;
	assign w3181 = w3182 ^ w3164;
	assign w3223 = w3229 ^ w3181;
	assign w3239 = w46124 ^ w3240;
	assign w3232 = w3241 & w3239;
	assign w3183 = w3226 ^ w3232;
	assign w3224 = w3183 ^ w3174;
	assign w3220 = w3224 & w3223;
	assign w3225 = w3247 & w3238;
	assign w43665 = w3225 ^ w3231;
	assign w3175 = w43665 ^ w3160;
	assign w3221 = w3183 ^ w3175;
	assign w3137 = w3169 ^ w43665;
	assign w3180 = w46119 ^ w3137;
	assign w3215 = w3220 ^ w3180;
	assign w3236 = w3166 ^ w3161;
	assign w3228 = w3243 & w3236;
	assign w43666 = w3225 ^ w3228;
	assign w3178 = w3226 ^ w43666;
	assign w3134 = w3229 ^ w3178;
	assign w3138 = w3164 ^ w43666;
	assign w3222 = w3138 ^ w3163;
	assign w3219 = w3220 ^ w3222;
	assign w3218 = w3221 & w3219;
	assign w3126 = w3218 ^ w3174;
	assign w3217 = w3218 ^ w3180;
	assign w3196 = w3217 & w3236;
	assign w3187 = w3217 & w3243;
	assign w3129 = w3218 ^ w3230;
	assign w3216 = w46123 ^ w3134;
	assign w3214 = w3215 & w3216;
	assign w3213 = w3214 ^ w3222;
	assign w3212 = w3220 ^ w3214;
	assign w3190 = w3213 & w3245;
	assign w3133 = w3214 ^ w3178;
	assign w3199 = w3213 & w46124;
	assign w3132 = w3214 ^ w3231;
	assign w3127 = w3132 ^ w3228;
	assign w3211 = w3222 & w3212;
	assign w3209 = w3211 ^ w3219;
	assign w43669 = w3211 ^ w3229;
	assign w3203 = w43669 ^ w3181;
	assign w3208 = w3217 & w3209;
	assign w3131 = w3208 ^ w3232;
	assign w3173 = w3208 ^ w3183;
	assign w3204 = w3173 ^ w3126;
	assign w3198 = w3204 & w3234;
	assign w3189 = w3204 & w3249;
	assign w3156 = w3198 ^ w3189;
	assign w3207 = w3173 ^ w3175;
	assign w3188 = w3207 & w3242;
	assign w3197 = w3207 & w3246;
	assign w3140 = w3196 ^ w3197;
	assign w43667 = w3197 ^ w3198;
	assign w3158 = w3196 ^ w3188;
	assign w3170 = w46123 ^ w43669;
	assign w3123 = w3170 ^ w3131;
	assign w3130 = w3160 ^ w3123;
	assign w3206 = w3127 ^ w3130;
	assign w3184 = w3206 & w3247;
	assign w3193 = w3206 & w3238;
	assign w3171 = w3189 ^ w3193;
	assign w3149 = ~w3171;
	assign w3148 = w3149 ^ w3187;
	assign w3125 = w3129 ^ w3165;
	assign w3128 = w46117 ^ w3125;
	assign w3124 = w46119 ^ w3125;
	assign w3202 = w3123 ^ w3124;
	assign w3194 = w3202 & w3235;
	assign w3179 = w3194 ^ w43667;
	assign w3155 = w3194 ^ w3197;
	assign w3152 = ~w3155;
	assign w3145 = w3190 ^ w3179;
	assign w3142 = ~w3145;
	assign w3205 = w3127 ^ w3128;
	assign w3195 = w3205 & w3237;
	assign w3150 = w3195 ^ w3184;
	assign w3146 = ~w3150;
	assign w3151 = w3194 ^ w3195;
	assign w3185 = w3202 & w3250;
	assign w3139 = w3195 ^ w3179;
	assign w3186 = w3205 & w3248;
	assign w43515 = w3185 ^ w3186;
	assign w3154 = w3158 ^ w43515;
	assign w3153 = w3149 ^ w3154;
	assign w3253 = w3152 ^ w3153;
	assign w46014 = ~w3253;
	assign w50963 = w46014 ^ w808;
	assign w3192 = w3203 & w3244;
	assign w3210 = w3170 ^ w3133;
	assign w3200 = w3210 & w3239;
	assign w3191 = w3210 & w3241;
	assign w3167 = w3191 ^ w43515;
	assign w3168 = w3192 ^ w3167;
	assign w46020 = w3168 ^ w3139;
	assign w50969 = w46020 ^ w814;
	assign w3172 = w3200 ^ w3168;
	assign w3141 = w3199 ^ w3172;
	assign w46016 = w3140 ^ w3141;
	assign w50965 = w46016 ^ w810;
	assign w3201 = w3203 & w3240;
	assign w43668 = w3199 ^ w3201;
	assign w3157 = w43668 ^ w3154;
	assign w3254 = w3156 ^ w3157;
	assign w46013 = ~w3254;
	assign w3144 = w3148 ^ w43668;
	assign w3147 = w3186 ^ w3144;
	assign w3251 = w3146 ^ w3147;
	assign w46018 = ~w3251;
	assign w50967 = w46018 ^ w812;
	assign w3177 = w3201 ^ w3172;
	assign w3252 = w3177 ^ w3151;
	assign w46019 = ~w3252;
	assign w46017 = w43667 ^ w3177;
	assign w50966 = w46017 ^ w811;
	assign w50968 = w46019 ^ w813;
	assign w3143 = w3167 ^ w3144;
	assign w46015 = w3142 ^ w3143;
	assign w50964 = w46015 ^ w809;
	assign w50962 = w46013 ^ w807;
	assign w10188 = w45851 ^ w45210;
	assign w10530 = w10187 ^ w10188;
	assign w50834 = w10530 ^ w10490;
	assign w46115 = w50834 ^ w624;
	assign w3383 = w46109 ^ w46115;
	assign w3293 = w46115 ^ w46113;
	assign w3374 = w3293 ^ w3382;
	assign w3373 = w46116 ^ w3374;
	assign w50839 = w45809 ^ w10403;
	assign w46110 = w50839 ^ w629;
	assign w3296 = w46112 ^ w46110;
	assign w3300 = w46116 ^ w46110;
	assign w3380 = w46111 ^ w3300;
	assign w3376 = w46115 ^ w3380;
	assign w3377 = w3294 ^ w3300;
	assign w3363 = w3380 & w3376;
	assign w3255 = w3296 ^ w46111;
	assign w3256 = w3296 ^ w3294;
	assign w3372 = w3293 ^ w3256;
	assign w3379 = w46116 ^ w3255;
	assign w3365 = w46116 & w3379;
	assign w45955 = ~w10435;
	assign w10398 = w45955 ^ w45850;
	assign w10426 = w45955 ^ w45809;
	assign w10395 = w45955 ^ w50906;
	assign w10393 = w10394 ^ w10395;
	assign w50844 = ~w10393;
	assign w50842 = w10397 ^ w10398;
	assign w46107 = w50842 ^ w632;
	assign w3510 = w46107 ^ w3514;
	assign w3444 = w46107 ^ w46106;
	assign w3512 = w3516 ^ w3444;
	assign w3509 = w3444 ^ w3511;
	assign w3497 = w3514 & w3510;
	assign w3517 = w46101 ^ w46107;
	assign w46105 = w50844 ^ w634;
	assign w3404 = w46105 ^ w46106;
	assign w3427 = w46107 ^ w46105;
	assign w3508 = w3427 ^ w3516;
	assign w3501 = w3508 & w3512;
	assign w3429 = w46106 ^ w3427;
	assign w3505 = w46102 ^ w3429;
	assign w3506 = w3427 ^ w3390;
	assign w3493 = w3515 & w3506;
	assign w3433 = w3501 ^ w3430;
	assign w3507 = w46108 ^ w3508;
	assign w3504 = w3434 ^ w3429;
	assign w3496 = w3511 & w3504;
	assign w43676 = w3493 ^ w3496;
	assign w3446 = w3494 ^ w43676;
	assign w3402 = w3497 ^ w3446;
	assign w3495 = w3516 & w3505;
	assign w3502 = w46103 ^ w3429;
	assign w3498 = w3517 & w3502;
	assign w3432 = w3498 ^ w3428;
	assign w3406 = w3432 ^ w43676;
	assign w3500 = w3509 & w3507;
	assign w50824 = w10426 ^ w10427;
	assign w46125 = w50824 ^ w614;
	assign w3115 = w46125 ^ w46131;
	assign w3113 = w46125 ^ w46130;
	assign w3114 = w46128 ^ w46125;
	assign w3106 = w3025 ^ w3114;
	assign w3105 = w46132 ^ w3106;
	assign w3026 = w46127 ^ w46125;
	assign w3101 = w3026 ^ w3116;
	assign w3109 = w3026 ^ w3032;
	assign w3107 = w3042 ^ w3109;
	assign w2988 = w3028 ^ w3026;
	assign w3104 = w3025 ^ w2988;
	assign w3091 = w3113 & w3104;
	assign w3110 = w3114 ^ w3042;
	assign w3099 = w3106 & w3110;
	assign w3031 = w3099 ^ w3028;
	assign w3093 = w3114 & w3103;
	assign w3029 = w3093 ^ w3027;
	assign w3035 = w3031 ^ w3029;
	assign w3040 = w46125 ^ w3035;
	assign w3098 = w3107 & w3105;
	assign w3094 = w3109 & w3102;
	assign w43659 = w3091 ^ w3094;
	assign w3096 = w3115 & w3100;
	assign w3030 = w3096 ^ w3026;
	assign w3004 = w3030 ^ w43659;
	assign w3088 = w3004 ^ w3029;
	assign w3484 = w46107 ^ w3402;
	assign w3431 = w3495 ^ w3429;
	assign w3490 = w3406 ^ w3431;
	assign w3092 = w3116 & w3101;
	assign w3044 = w3092 ^ w43659;
	assign w3000 = w3095 ^ w3044;
	assign w3049 = w3092 ^ w3098;
	assign w3001 = w3092 ^ w3093;
	assign w3048 = w3001 ^ w3002;
	assign w3047 = w3048 ^ w3030;
	assign w3089 = w3095 ^ w3047;
	assign w3090 = w3049 ^ w3040;
	assign w3086 = w3090 & w3089;
	assign w3082 = w46131 ^ w3000;
	assign w43679 = w3493 ^ w3499;
	assign w3443 = w43679 ^ w3428;
	assign w3437 = w3433 ^ w3431;
	assign w3405 = w3437 ^ w43679;
	assign w3448 = w46103 ^ w3405;
	assign w3442 = w46101 ^ w3437;
	assign w3451 = w3494 ^ w3500;
	assign w3492 = w3451 ^ w3442;
	assign w3489 = w3451 ^ w3443;
	assign w3403 = w3494 ^ w3495;
	assign w3450 = w3403 ^ w3404;
	assign w3449 = w3450 ^ w3432;
	assign w3491 = w3497 ^ w3449;
	assign w3488 = w3492 & w3491;
	assign w3483 = w3488 ^ w3448;
	assign w3482 = w3483 & w3484;
	assign w3480 = w3488 ^ w3482;
	assign w3487 = w3488 ^ w3490;
	assign w3479 = w3490 & w3480;
	assign w3477 = w3479 ^ w3487;
	assign w43678 = w3479 ^ w3497;
	assign w3400 = w3482 ^ w3499;
	assign w3395 = w3400 ^ w3496;
	assign w3486 = w3489 & w3487;
	assign w3485 = w3486 ^ w3448;
	assign w3476 = w3485 & w3477;
	assign w3455 = w3485 & w3511;
	assign w3399 = w3476 ^ w3500;
	assign w3441 = w3476 ^ w3451;
	assign w3397 = w3486 ^ w3498;
	assign w3393 = w3397 ^ w3433;
	assign w3392 = w46103 ^ w3393;
	assign w3396 = w46101 ^ w3393;
	assign w3473 = w3395 ^ w3396;
	assign w3394 = w3486 ^ w3442;
	assign w3472 = w3441 ^ w3394;
	assign w3466 = w3472 & w3502;
	assign w3457 = w3472 & w3517;
	assign w3424 = w3466 ^ w3457;
	assign w3438 = w46107 ^ w43678;
	assign w3391 = w3438 ^ w3399;
	assign w3470 = w3391 ^ w3392;
	assign w3462 = w3470 & w3503;
	assign w3471 = w43678 ^ w3449;
	assign w3469 = w3471 & w3508;
	assign w3464 = w3485 & w3504;
	assign w3398 = w3428 ^ w3391;
	assign w3481 = w3482 ^ w3490;
	assign w3467 = w3481 & w46108;
	assign w3458 = w3481 & w3513;
	assign w43681 = w3467 ^ w3469;
	assign w3463 = w3473 & w3505;
	assign w3419 = w3462 ^ w3463;
	assign w3453 = w3470 & w3518;
	assign w3475 = w3441 ^ w3443;
	assign w3465 = w3475 & w3514;
	assign w3408 = w3464 ^ w3465;
	assign w3423 = w3462 ^ w3465;
	assign w3456 = w3475 & w3510;
	assign w3426 = w3464 ^ w3456;
	assign w3420 = ~w3423;
	assign w43680 = w3465 ^ w3466;
	assign w3447 = w3462 ^ w43680;
	assign w3413 = w3458 ^ w3447;
	assign w3410 = ~w3413;
	assign w3454 = w3473 & w3516;
	assign w43677 = w3453 ^ w3454;
	assign w3422 = w3426 ^ w43677;
	assign w3425 = w43681 ^ w3422;
	assign w3401 = w3482 ^ w3446;
	assign w3478 = w3438 ^ w3401;
	assign w3468 = w3478 & w3507;
	assign w3459 = w3478 & w3509;
	assign w3435 = w3459 ^ w43677;
	assign w3407 = w3463 ^ w3447;
	assign w3085 = w3086 ^ w3088;
	assign w3522 = w3424 ^ w3425;
	assign w46093 = ~w3522;
	assign w51042 = w46093 ^ w759;
	assign w3474 = w3395 ^ w3398;
	assign w3461 = w3474 & w3506;
	assign w3452 = w3474 & w3515;
	assign w3418 = w3463 ^ w3452;
	assign w3439 = w3457 ^ w3461;
	assign w3417 = ~w3439;
	assign w3421 = w3417 ^ w3422;
	assign w3521 = w3420 ^ w3421;
	assign w3416 = w3417 ^ w3455;
	assign w3412 = w3416 ^ w43681;
	assign w3411 = w3435 ^ w3412;
	assign w46095 = w3410 ^ w3411;
	assign w51044 = w46095 ^ w761;
	assign w46094 = ~w3521;
	assign w3415 = w3454 ^ w3412;
	assign w3414 = ~w3418;
	assign w3519 = w3414 ^ w3415;
	assign w46098 = ~w3519;
	assign w51047 = w46098 ^ w764;
	assign w51043 = w46094 ^ w760;
	assign w43662 = w3091 ^ w3097;
	assign w3003 = w3035 ^ w43662;
	assign w3046 = w46127 ^ w3003;
	assign w3081 = w3086 ^ w3046;
	assign w3080 = w3081 & w3082;
	assign w3079 = w3080 ^ w3088;
	assign w3056 = w3079 & w3111;
	assign w3065 = w3079 & w46132;
	assign w3078 = w3086 ^ w3080;
	assign w2998 = w3080 ^ w3097;
	assign w2993 = w2998 ^ w3094;
	assign w3077 = w3088 & w3078;
	assign w43661 = w3077 ^ w3095;
	assign w3036 = w46131 ^ w43661;
	assign w3075 = w3077 ^ w3085;
	assign w2999 = w3080 ^ w3044;
	assign w3076 = w3036 ^ w2999;
	assign w3057 = w3076 & w3107;
	assign w3066 = w3076 & w3105;
	assign w3069 = w43661 ^ w3047;
	assign w3067 = w3069 & w3106;
	assign w43664 = w3065 ^ w3067;
	assign w3058 = w3069 & w3110;
	assign w3041 = w43662 ^ w3026;
	assign w3087 = w3049 ^ w3041;
	assign w3084 = w3087 & w3085;
	assign w3083 = w3084 ^ w3046;
	assign w3053 = w3083 & w3109;
	assign w2992 = w3084 ^ w3040;
	assign w3062 = w3083 & w3102;
	assign w3074 = w3083 & w3075;
	assign w3039 = w3074 ^ w3049;
	assign w3070 = w3039 ^ w2992;
	assign w3064 = w3070 & w3100;
	assign w3073 = w3039 ^ w3041;
	assign w3055 = w3070 & w3115;
	assign w3022 = w3064 ^ w3055;
	assign w2995 = w3084 ^ w3096;
	assign w2991 = w2995 ^ w3031;
	assign w2994 = w46125 ^ w2991;
	assign w3071 = w2993 ^ w2994;
	assign w2990 = w46127 ^ w2991;
	assign w3052 = w3071 & w3114;
	assign w3061 = w3071 & w3103;
	assign w3054 = w3073 & w3108;
	assign w3024 = w3062 ^ w3054;
	assign w3063 = w3073 & w3112;
	assign w3006 = w3062 ^ w3063;
	assign w2997 = w3074 ^ w3098;
	assign w2989 = w3036 ^ w2997;
	assign w2996 = w3026 ^ w2989;
	assign w3068 = w2989 ^ w2990;
	assign w3060 = w3068 & w3101;
	assign w3017 = w3060 ^ w3061;
	assign w3051 = w3068 & w3116;
	assign w3021 = w3060 ^ w3063;
	assign w43660 = w3051 ^ w3052;
	assign w3033 = w3057 ^ w43660;
	assign w3020 = w3024 ^ w43660;
	assign w3018 = ~w3021;
	assign w3072 = w2993 ^ w2996;
	assign w3050 = w3072 & w3113;
	assign w3016 = w3061 ^ w3050;
	assign w3012 = ~w3016;
	assign w3059 = w3072 & w3104;
	assign w3037 = w3055 ^ w3059;
	assign w3015 = ~w3037;
	assign w3019 = w3015 ^ w3020;
	assign w3014 = w3015 ^ w3053;
	assign w3119 = w3018 ^ w3019;
	assign w46038 = ~w3119;
	assign w3010 = w3014 ^ w43664;
	assign w3009 = w3033 ^ w3010;
	assign w3013 = w3052 ^ w3010;
	assign w3117 = w3012 ^ w3013;
	assign w46042 = ~w3117;
	assign w50991 = w46042 ^ w772;
	assign w3023 = w43664 ^ w3020;
	assign w3120 = w3022 ^ w3023;
	assign w46037 = ~w3120;
	assign w50986 = w46037 ^ w767;
	assign w50987 = w46038 ^ w768;
	assign w3034 = w3058 ^ w3033;
	assign w3038 = w3066 ^ w3034;
	assign w3007 = w3065 ^ w3038;
	assign w3043 = w3067 ^ w3038;
	assign w46040 = w3006 ^ w3007;
	assign w3118 = w3043 ^ w3017;
	assign w46043 = ~w3118;
	assign w50992 = w46043 ^ w773;
	assign w50989 = w46040 ^ w770;
	assign w43663 = w3063 ^ w3064;
	assign w46041 = w43663 ^ w3043;
	assign w50990 = w46041 ^ w771;
	assign w3045 = w3060 ^ w43663;
	assign w3005 = w3061 ^ w3045;
	assign w3011 = w3056 ^ w3045;
	assign w3008 = ~w3011;
	assign w46039 = w3008 ^ w3009;
	assign w50988 = w46039 ^ w769;
	assign w46044 = w3034 ^ w3005;
	assign w50993 = w46044 ^ w774;
	assign w45960 = ~w10442;
	assign w10387 = w45960 ^ w50851;
	assign w10366 = w45960 ^ w50868;
	assign w50744 = w10366 ^ w10367;
	assign w46205 = w50744 ^ w726;
	assign w2445 = w46205 ^ w46211;
	assign w2426 = w2445 & w2430;
	assign w10230 = w45960 ^ w45845;
	assign w10512 = w10230 ^ w10231;
	assign w2356 = w46207 ^ w46205;
	assign w2360 = w2426 ^ w2356;
	assign w2318 = w2358 ^ w2356;
	assign w2431 = w2356 ^ w2446;
	assign w2422 = w2446 & w2431;
	assign w2443 = w46205 ^ w46210;
	assign w2439 = w2356 ^ w2362;
	assign w2437 = w2372 ^ w2439;
	assign w2424 = w2439 & w2432;
	assign w2444 = w46208 ^ w46205;
	assign w2423 = w2444 & w2433;
	assign w2440 = w2444 ^ w2372;
	assign w2331 = w2422 ^ w2423;
	assign w2378 = w2331 ^ w2332;
	assign w2377 = w2378 ^ w2360;
	assign w2419 = w2425 ^ w2377;
	assign w2359 = w2423 ^ w2357;
	assign w50730 = w10512 ^ w10504;
	assign w46219 = w50730 ^ w712;
	assign w2221 = w46219 ^ w46217;
	assign w2223 = w46218 ^ w2221;
	assign w2298 = w2228 ^ w2223;
	assign w2299 = w46214 ^ w2223;
	assign w2296 = w46215 ^ w2223;
	assign w2238 = w46219 ^ w46218;
	assign w2303 = w2238 ^ w2305;
	assign w2290 = w2305 & w2298;
	assign w2311 = w46213 ^ w46219;
	assign w2292 = w2311 & w2296;
	assign w2226 = w2292 ^ w2222;
	assign w2434 = w2355 ^ w2318;
	assign w2421 = w2443 & w2434;
	assign w43632 = w2421 ^ w2424;
	assign w2334 = w2360 ^ w43632;
	assign w43631 = w2421 ^ w2427;
	assign w2374 = w2422 ^ w43632;
	assign w2330 = w2425 ^ w2374;
	assign w2412 = w46211 ^ w2330;
	assign w2304 = w46219 ^ w2308;
	assign w2291 = w2308 & w2304;
	assign w2371 = w43631 ^ w2356;
	assign w2436 = w2355 ^ w2444;
	assign w2435 = w46212 ^ w2436;
	assign w2428 = w2437 & w2435;
	assign w2379 = w2422 ^ w2428;
	assign w2417 = w2379 ^ w2371;
	assign w2429 = w2436 & w2440;
	assign w2361 = w2429 ^ w2358;
	assign w2365 = w2361 ^ w2359;
	assign w2370 = w46205 ^ w2365;
	assign w2420 = w2379 ^ w2370;
	assign w2416 = w2420 & w2419;
	assign w2333 = w2365 ^ w43631;
	assign w2376 = w46207 ^ w2333;
	assign w2411 = w2416 ^ w2376;
	assign w2410 = w2411 & w2412;
	assign w2328 = w2410 ^ w2427;
	assign w2408 = w2416 ^ w2410;
	assign w2323 = w2328 ^ w2424;
	assign w2329 = w2410 ^ w2374;
	assign w2418 = w2334 ^ w2359;
	assign w2409 = w2410 ^ w2418;
	assign w2386 = w2409 & w2441;
	assign w2407 = w2418 & w2408;
	assign w2415 = w2416 ^ w2418;
	assign w2405 = w2407 ^ w2415;
	assign w2395 = w2409 & w46212;
	assign w43635 = w2407 ^ w2425;
	assign w2399 = w43635 ^ w2377;
	assign w2388 = w2399 & w2440;
	assign w2397 = w2399 & w2436;
	assign w2366 = w46211 ^ w43635;
	assign w2406 = w2366 ^ w2329;
	assign w2387 = w2406 & w2437;
	assign w2396 = w2406 & w2435;
	assign w2414 = w2417 & w2415;
	assign w2325 = w2414 ^ w2426;
	assign w2322 = w2414 ^ w2370;
	assign w2413 = w2414 ^ w2376;
	assign w2404 = w2413 & w2405;
	assign w2327 = w2404 ^ w2428;
	assign w2319 = w2366 ^ w2327;
	assign w2326 = w2356 ^ w2319;
	assign w2402 = w2323 ^ w2326;
	assign w2369 = w2404 ^ w2379;
	assign w2403 = w2369 ^ w2371;
	assign w2384 = w2403 & w2438;
	assign w2400 = w2369 ^ w2322;
	assign w2392 = w2413 & w2432;
	assign w2380 = w2402 & w2443;
	assign w2385 = w2400 & w2445;
	assign w2393 = w2403 & w2442;
	assign w2383 = w2413 & w2439;
	assign w2354 = w2392 ^ w2384;
	assign w2394 = w2400 & w2430;
	assign w43633 = w2393 ^ w2394;
	assign w43634 = w2395 ^ w2397;
	assign w2336 = w2392 ^ w2393;
	assign w2321 = w2325 ^ w2361;
	assign w2320 = w46207 ^ w2321;
	assign w2398 = w2319 ^ w2320;
	assign w2381 = w2398 & w2446;
	assign w2390 = w2398 & w2431;
	assign w2375 = w2390 ^ w43633;
	assign w2341 = w2386 ^ w2375;
	assign w2351 = w2390 ^ w2393;
	assign w2348 = ~w2351;
	assign w2338 = ~w2341;
	assign w2324 = w46205 ^ w2321;
	assign w2401 = w2323 ^ w2324;
	assign w2391 = w2401 & w2433;
	assign w2346 = w2391 ^ w2380;
	assign w2347 = w2390 ^ w2391;
	assign w2382 = w2401 & w2444;
	assign w43513 = w2381 ^ w2382;
	assign w2350 = w2354 ^ w43513;
	assign w2353 = w43634 ^ w2350;
	assign w2335 = w2391 ^ w2375;
	assign w2342 = ~w2346;
	assign w2363 = w2387 ^ w43513;
	assign w2364 = w2388 ^ w2363;
	assign w46028 = w2364 ^ w2335;
	assign w50977 = w46028 ^ w822;
	assign w2368 = w2396 ^ w2364;
	assign w2373 = w2397 ^ w2368;
	assign w2448 = w2373 ^ w2347;
	assign w46027 = ~w2448;
	assign w46025 = w43633 ^ w2373;
	assign w50974 = w46025 ^ w819;
	assign w50976 = w46027 ^ w821;
	assign w2337 = w2395 ^ w2368;
	assign w46024 = w2336 ^ w2337;
	assign w50973 = w46024 ^ w818;
	assign w2389 = w2402 & w2434;
	assign w2367 = w2385 ^ w2389;
	assign w2345 = ~w2367;
	assign w2344 = w2345 ^ w2383;
	assign w2349 = w2345 ^ w2350;
	assign w2449 = w2348 ^ w2349;
	assign w46022 = ~w2449;
	assign w50971 = w46022 ^ w816;
	assign w2340 = w2344 ^ w43634;
	assign w2339 = w2363 ^ w2340;
	assign w46023 = w2338 ^ w2339;
	assign w2343 = w2382 ^ w2340;
	assign w50972 = w46023 ^ w817;
	assign w2447 = w2342 ^ w2343;
	assign w46026 = ~w2447;
	assign w50975 = w46026 ^ w820;
	assign w2352 = w2394 ^ w2385;
	assign w2450 = w2352 ^ w2353;
	assign w46021 = ~w2450;
	assign w50970 = w46021 ^ w815;
	assign w50733 = w10386 ^ w10387;
	assign w46216 = w50733 ^ w715;
	assign w2312 = w46218 ^ w46216;
	assign w2224 = w46216 ^ w46214;
	assign w2184 = w2224 ^ w2222;
	assign w2183 = w2224 ^ w46215;
	assign w2307 = w46220 ^ w2183;
	assign w2293 = w46220 & w2307;
	assign w2300 = w2221 ^ w2184;
	assign w2287 = w2309 & w2300;
	assign w43625 = w2287 ^ w2290;
	assign w43628 = w2287 ^ w2293;
	assign w2200 = w2226 ^ w43625;
	assign w2297 = w2222 ^ w2312;
	assign w2288 = w2312 & w2297;
	assign w2240 = w2288 ^ w43625;
	assign w2196 = w2291 ^ w2240;
	assign w2278 = w46219 ^ w2196;
	assign w2237 = w43628 ^ w2222;
	assign w2310 = w46216 ^ w46213;
	assign w2289 = w2310 & w2299;
	assign w2197 = w2288 ^ w2289;
	assign w2244 = w2197 ^ w2198;
	assign w2243 = w2244 ^ w2226;
	assign w2306 = w2310 ^ w2238;
	assign w2302 = w2221 ^ w2310;
	assign w2225 = w2289 ^ w2223;
	assign w2284 = w2200 ^ w2225;
	assign w2295 = w2302 & w2306;
	assign w2227 = w2295 ^ w2224;
	assign w2231 = w2227 ^ w2225;
	assign w2199 = w2231 ^ w43628;
	assign w2236 = w46213 ^ w2231;
	assign w2242 = w46215 ^ w2199;
	assign w2301 = w46220 ^ w2302;
	assign w2294 = w2303 & w2301;
	assign w2285 = w2291 ^ w2243;
	assign w2245 = w2288 ^ w2294;
	assign w2286 = w2245 ^ w2236;
	assign w2282 = w2286 & w2285;
	assign w2281 = w2282 ^ w2284;
	assign w2277 = w2282 ^ w2242;
	assign w2276 = w2277 & w2278;
	assign w2274 = w2282 ^ w2276;
	assign w2273 = w2284 & w2274;
	assign w43627 = w2273 ^ w2291;
	assign w2232 = w46219 ^ w43627;
	assign w2265 = w43627 ^ w2243;
	assign w2263 = w2265 & w2302;
	assign w2254 = w2265 & w2306;
	assign w2275 = w2276 ^ w2284;
	assign w2252 = w2275 & w2307;
	assign w2261 = w2275 & w46220;
	assign w2195 = w2276 ^ w2240;
	assign w2272 = w2232 ^ w2195;
	assign w2253 = w2272 & w2303;
	assign w2262 = w2272 & w2301;
	assign w43630 = w2261 ^ w2263;
	assign w2271 = w2273 ^ w2281;
	assign w2194 = w2276 ^ w2293;
	assign w2189 = w2194 ^ w2290;
	assign w2283 = w2245 ^ w2237;
	assign w2280 = w2281 & w2283;
	assign w2188 = w2280 ^ w2236;
	assign w2191 = w2280 ^ w2292;
	assign w2279 = w2280 ^ w2242;
	assign w2258 = w2279 & w2298;
	assign w2270 = w2279 & w2271;
	assign w2193 = w2270 ^ w2294;
	assign w2235 = w2270 ^ w2245;
	assign w2269 = w2235 ^ w2237;
	assign w2250 = w2269 & w2304;
	assign w2220 = w2258 ^ w2250;
	assign w2266 = w2235 ^ w2188;
	assign w2185 = w2232 ^ w2193;
	assign w2260 = w2266 & w2296;
	assign w2251 = w2266 & w2311;
	assign w2218 = w2260 ^ w2251;
	assign w2249 = w2279 & w2305;
	assign w2192 = w2222 ^ w2185;
	assign w2268 = w2189 ^ w2192;
	assign w2246 = w2268 & w2309;
	assign w2255 = w2268 & w2300;
	assign w2233 = w2251 ^ w2255;
	assign w2211 = ~w2233;
	assign w2210 = w2211 ^ w2249;
	assign w2206 = w2210 ^ w43630;
	assign w2259 = w2269 & w2308;
	assign w43629 = w2259 ^ w2260;
	assign w2202 = w2258 ^ w2259;
	assign w2187 = w2191 ^ w2227;
	assign w2186 = w46215 ^ w2187;
	assign w2264 = w2185 ^ w2186;
	assign w2247 = w2264 & w2312;
	assign w2190 = w46213 ^ w2187;
	assign w2267 = w2189 ^ w2190;
	assign w2257 = w2267 & w2299;
	assign w2212 = w2257 ^ w2246;
	assign w2208 = ~w2212;
	assign w2248 = w2267 & w2310;
	assign w43626 = w2247 ^ w2248;
	assign w2209 = w2248 ^ w2206;
	assign w2313 = w2208 ^ w2209;
	assign w2229 = w2253 ^ w43626;
	assign w2205 = w2229 ^ w2206;
	assign w46050 = ~w2313;
	assign w50999 = w46050 ^ w780;
	assign w2230 = w2254 ^ w2229;
	assign w2234 = w2262 ^ w2230;
	assign w2203 = w2261 ^ w2234;
	assign w46048 = w2202 ^ w2203;
	assign w50997 = w46048 ^ w778;
	assign w2239 = w2263 ^ w2234;
	assign w46049 = w43629 ^ w2239;
	assign w50998 = w46049 ^ w779;
	assign w2216 = w2220 ^ w43626;
	assign w2219 = w43630 ^ w2216;
	assign w2316 = w2218 ^ w2219;
	assign w46045 = ~w2316;
	assign w50994 = w46045 ^ w775;
	assign w2215 = w2211 ^ w2216;
	assign w39809 = w39839 & w39865;
	assign w39770 = w39771 ^ w39809;
	assign w39766 = w39770 ^ w45043;
	assign w39765 = w39789 ^ w39766;
	assign w50901 = w39764 ^ w39765;
	assign w10269 = w10271 ^ w50901;
	assign w50803 = w10269 ^ w10270;
	assign w46146 = w50803 ^ w657;
	assign w40408 = w46146 ^ w46144;
	assign w40319 = w46146 ^ w40317;
	assign w40394 = w40324 ^ w40319;
	assign w40294 = w46145 ^ w46146;
	assign w40334 = w46147 ^ w46146;
	assign w40402 = w40406 ^ w40334;
	assign w40391 = w40398 & w40402;
	assign w40323 = w40391 ^ w40320;
	assign w40395 = w46142 ^ w40319;
	assign w40385 = w40406 & w40395;
	assign w40321 = w40385 ^ w40319;
	assign w10215 = w10214 ^ w50901;
	assign w10518 = w10215 ^ w10216;
	assign w50788 = w10518 ^ w10477;
	assign w46161 = w50788 ^ w642;
	assign w42059 = w46163 ^ w46161;
	assign w42140 = w42059 ^ w42148;
	assign w40405 = w46141 ^ w46146;
	assign w40327 = w40323 ^ w40321;
	assign w40332 = w46141 ^ w40327;
	assign w10487 = w50897 ^ w50901;
	assign w10300 = ~w10487;
	assign w10298 = w10300 ^ w45823;
	assign w50787 = w10298 ^ w10299;
	assign w46162 = w50787 ^ w641;
	assign w42076 = w46163 ^ w46162;
	assign w42144 = w42148 ^ w42076;
	assign w42147 = w46157 ^ w46162;
	assign w42133 = w42140 & w42144;
	assign w42061 = w46162 ^ w42059;
	assign w42150 = w46162 ^ w46160;
	assign w10282 = w10502 ^ w10487;
	assign w50795 = w50886 ^ w10282;
	assign w46154 = w50795 ^ w649;
	assign w40964 = w46153 ^ w46154;
	assign w41004 = w46155 ^ w46154;
	assign w41072 = w41076 ^ w41004;
	assign w41061 = w41068 & w41072;
	assign w40993 = w41061 ^ w40990;
	assign w41075 = w46149 ^ w46154;
	assign w40989 = w46154 ^ w40987;
	assign w41065 = w46150 ^ w40989;
	assign w41064 = w40994 ^ w40989;
	assign w41055 = w41076 & w41065;
	assign w40991 = w41055 ^ w40989;
	assign w40997 = w40993 ^ w40991;
	assign w41002 = w46149 ^ w40997;
	assign w41078 = w46154 ^ w46152;
	assign w42036 = w46161 ^ w46162;
	assign w10253 = w10255 ^ w10487;
	assign w50812 = w10253 ^ w10254;
	assign w46137 = w50812 ^ w666;
	assign w39647 = w46139 ^ w46137;
	assign w39624 = w46137 ^ w46138;
	assign w39728 = w39647 ^ w39736;
	assign w39649 = w46138 ^ w39647;
	assign w39722 = w46135 ^ w39649;
	assign w39727 = w46140 ^ w39728;
	assign w39718 = w39737 & w39722;
	assign w39652 = w39718 ^ w39648;
	assign w39721 = w39728 & w39732;
	assign w39769 = w39808 ^ w39766;
	assign w39873 = w39768 ^ w39769;
	assign w45829 = ~w39873;
	assign w10462 = w45860 ^ w45829;
	assign w10297 = w10462 ^ w50903;
	assign w10295 = ~w10297;
	assign w50790 = w10295 ^ w10296;
	assign w46159 = w50790 ^ w644;
	assign w10290 = w10451 ^ w45829;
	assign w10289 = w10290 ^ w10291;
	assign w50791 = ~w10289;
	assign w46158 = w50791 ^ w645;
	assign w42137 = w46158 ^ w42061;
	assign w42066 = w46164 ^ w46158;
	assign w10248 = w10466 ^ w10462;
	assign w42060 = w46159 ^ w46157;
	assign w42143 = w42060 ^ w42066;
	assign w42141 = w42076 ^ w42143;
	assign w10267 = w10473 ^ w45829;
	assign w50806 = w10267 ^ w10268;
	assign w46143 = w50806 ^ w660;
	assign w40279 = w40320 ^ w46143;
	assign w40404 = w46143 ^ w40324;
	assign w40403 = w46148 ^ w40279;
	assign w40389 = w46148 & w40403;
	assign w40318 = w46143 ^ w46141;
	assign w40280 = w40320 ^ w40318;
	assign w40396 = w40317 ^ w40280;
	assign w40401 = w40318 ^ w40324;
	assign w40399 = w40334 ^ w40401;
	assign w40386 = w40401 & w40394;
	assign w42127 = w42148 & w42137;
	assign w42063 = w42127 ^ w42061;
	assign w40400 = w46147 ^ w40404;
	assign w40387 = w40404 & w40400;
	assign w42062 = w46160 ^ w46158;
	assign w42021 = w42062 ^ w46159;
	assign w42145 = w46164 ^ w42021;
	assign w42131 = w46164 & w42145;
	assign w42022 = w42062 ^ w42060;
	assign w42138 = w42059 ^ w42022;
	assign w42125 = w42147 & w42138;
	assign w45136 = w42125 ^ w42131;
	assign w42075 = w45136 ^ w42060;
	assign w42136 = w42066 ^ w42061;
	assign w10277 = w10480 ^ w10462;
	assign w50798 = w45852 ^ w10277;
	assign w46151 = w50798 ^ w652;
	assign w40988 = w46151 ^ w46149;
	assign w41063 = w40988 ^ w41078;
	assign w41071 = w40988 ^ w40994;
	assign w41056 = w41071 & w41064;
	assign w41074 = w46151 ^ w40994;
	assign w41070 = w46155 ^ w41074;
	assign w41057 = w41074 & w41070;
	assign w41062 = w46151 ^ w40989;
	assign w40950 = w40990 ^ w40988;
	assign w41066 = w40987 ^ w40950;
	assign w41053 = w41075 & w41066;
	assign w45090 = w41053 ^ w41056;
	assign w41054 = w41078 & w41063;
	assign w40963 = w41054 ^ w41055;
	assign w41058 = w41077 & w41062;
	assign w41010 = w40963 ^ w40964;
	assign w41006 = w41054 ^ w45090;
	assign w40962 = w41057 ^ w41006;
	assign w40992 = w41058 ^ w40988;
	assign w40966 = w40992 ^ w45090;
	assign w41050 = w40966 ^ w40991;
	assign w41009 = w41010 ^ w40992;
	assign w40393 = w40318 ^ w40408;
	assign w40384 = w40408 & w40393;
	assign w40293 = w40384 ^ w40385;
	assign w40340 = w40293 ^ w40294;
	assign w40392 = w46143 ^ w40319;
	assign w40388 = w40407 & w40392;
	assign w40322 = w40388 ^ w40318;
	assign w40339 = w40340 ^ w40322;
	assign w40381 = w40387 ^ w40339;
	assign w41069 = w41004 ^ w41071;
	assign w41060 = w41069 & w41067;
	assign w41044 = w46155 ^ w40962;
	assign w41051 = w41057 ^ w41009;
	assign w42065 = w42133 ^ w42062;
	assign w42069 = w42065 ^ w42063;
	assign w42037 = w42069 ^ w45136;
	assign w42080 = w46159 ^ w42037;
	assign w40949 = w40990 ^ w46151;
	assign w41073 = w46156 ^ w40949;
	assign w41059 = w46156 & w41073;
	assign w45089 = w41053 ^ w41059;
	assign w40965 = w40997 ^ w45089;
	assign w41008 = w46151 ^ w40965;
	assign w42074 = w46157 ^ w42069;
	assign w40383 = w40405 & w40396;
	assign w45062 = w40383 ^ w40386;
	assign w40296 = w40322 ^ w45062;
	assign w40336 = w40384 ^ w45062;
	assign w40292 = w40387 ^ w40336;
	assign w40374 = w46147 ^ w40292;
	assign w40380 = w40296 ^ w40321;
	assign w42134 = w46159 ^ w42061;
	assign w42130 = w42149 & w42134;
	assign w42064 = w42130 ^ w42060;
	assign w41011 = w41054 ^ w41060;
	assign w41052 = w41011 ^ w41002;
	assign w41048 = w41052 & w41051;
	assign w41047 = w41048 ^ w41050;
	assign w41043 = w41048 ^ w41008;
	assign w41042 = w41043 & w41044;
	assign w40961 = w41042 ^ w41006;
	assign w41041 = w41042 ^ w41050;
	assign w41018 = w41041 & w41073;
	assign w41027 = w41041 & w46156;
	assign w40960 = w41042 ^ w41059;
	assign w40955 = w40960 ^ w41056;
	assign w41040 = w41048 ^ w41042;
	assign w41039 = w41050 & w41040;
	assign w45093 = w41039 ^ w41057;
	assign w41031 = w45093 ^ w41009;
	assign w41020 = w41031 & w41072;
	assign w40998 = w46155 ^ w45093;
	assign w41037 = w41039 ^ w41047;
	assign w41029 = w41031 & w41068;
	assign w45092 = w41027 ^ w41029;
	assign w42128 = w42143 & w42136;
	assign w45133 = w42125 ^ w42128;
	assign w42038 = w42064 ^ w45133;
	assign w42122 = w42038 ^ w42063;
	assign w41003 = w45089 ^ w40988;
	assign w41049 = w41011 ^ w41003;
	assign w41046 = w41049 & w41047;
	assign w40954 = w41046 ^ w41002;
	assign w41045 = w41046 ^ w41008;
	assign w41024 = w41045 & w41064;
	assign w41036 = w41045 & w41037;
	assign w41001 = w41036 ^ w41011;
	assign w41032 = w41001 ^ w40954;
	assign w41017 = w41032 & w41077;
	assign w41035 = w41001 ^ w41003;
	assign w41025 = w41035 & w41074;
	assign w41015 = w41045 & w41071;
	assign w41026 = w41032 & w41062;
	assign w45091 = w41025 ^ w41026;
	assign w40984 = w41026 ^ w41017;
	assign w41016 = w41035 & w41070;
	assign w40986 = w41024 ^ w41016;
	assign w40959 = w41036 ^ w41060;
	assign w40968 = w41024 ^ w41025;
	assign w40957 = w41046 ^ w41058;
	assign w40953 = w40957 ^ w40993;
	assign w40956 = w46149 ^ w40953;
	assign w40952 = w46151 ^ w40953;
	assign w41033 = w40955 ^ w40956;
	assign w41014 = w41033 & w41076;
	assign w41023 = w41033 & w41065;
	assign w50815 = w45861 ^ w10248;
	assign w46134 = w50815 ^ w669;
	assign w39650 = w46136 ^ w46134;
	assign w39653 = w39721 ^ w39650;
	assign w39654 = w46140 ^ w46134;
	assign w39734 = w46135 ^ w39654;
	assign w39730 = w46139 ^ w39734;
	assign w39731 = w39648 ^ w39654;
	assign w39729 = w39664 ^ w39731;
	assign w39720 = w39729 & w39727;
	assign w39717 = w39734 & w39730;
	assign w39671 = w39714 ^ w39720;
	assign w39609 = w39650 ^ w46135;
	assign w39733 = w46140 ^ w39609;
	assign w39610 = w39650 ^ w39648;
	assign w39726 = w39647 ^ w39610;
	assign w39713 = w39735 & w39726;
	assign w39725 = w46134 ^ w39649;
	assign w39715 = w39736 & w39725;
	assign w39623 = w39714 ^ w39715;
	assign w39670 = w39623 ^ w39624;
	assign w39651 = w39715 ^ w39649;
	assign w39657 = w39653 ^ w39651;
	assign w39662 = w46133 ^ w39657;
	assign w39719 = w46140 & w39733;
	assign w45032 = w39713 ^ w39719;
	assign w39663 = w45032 ^ w39648;
	assign w39709 = w39671 ^ w39663;
	assign w39625 = w39657 ^ w45032;
	assign w39668 = w46135 ^ w39625;
	assign w39669 = w39670 ^ w39652;
	assign w39711 = w39717 ^ w39669;
	assign w41038 = w40998 ^ w40961;
	assign w41019 = w41038 & w41069;
	assign w41028 = w41038 & w41067;
	assign w40951 = w40998 ^ w40959;
	assign w41030 = w40951 ^ w40952;
	assign w41022 = w41030 & w41063;
	assign w40983 = w41022 ^ w41025;
	assign w40979 = w41022 ^ w41023;
	assign w41013 = w41030 & w41078;
	assign w41007 = w41022 ^ w45091;
	assign w40967 = w41023 ^ w41007;
	assign w40973 = w41018 ^ w41007;
	assign w40970 = ~w40973;
	assign w43612 = w41013 ^ w41014;
	assign w40982 = w40986 ^ w43612;
	assign w40985 = w45092 ^ w40982;
	assign w41082 = w40984 ^ w40985;
	assign w40958 = w40988 ^ w40951;
	assign w41034 = w40955 ^ w40958;
	assign w41021 = w41034 & w41066;
	assign w41012 = w41034 & w41075;
	assign w40978 = w41023 ^ w41012;
	assign w40974 = ~w40978;
	assign w45981 = ~w41082;
	assign w50930 = w45981 ^ w839;
	assign w40995 = w41019 ^ w43612;
	assign w40996 = w41020 ^ w40995;
	assign w41000 = w41028 ^ w40996;
	assign w41005 = w41029 ^ w41000;
	assign w40969 = w41027 ^ w41000;
	assign w45985 = w45091 ^ w41005;
	assign w50934 = w45985 ^ w843;
	assign w41080 = w41005 ^ w40979;
	assign w45987 = ~w41080;
	assign w50936 = w45987 ^ w845;
	assign w45984 = w40968 ^ w40969;
	assign w50933 = w45984 ^ w842;
	assign w40980 = ~w40983;
	assign w45988 = w40996 ^ w40967;
	assign w50937 = w45988 ^ w846;
	assign w40999 = w41017 ^ w41021;
	assign w40977 = ~w40999;
	assign w40981 = w40977 ^ w40982;
	assign w41081 = w40980 ^ w40981;
	assign w45982 = ~w41081;
	assign w50931 = w45982 ^ w840;
	assign w40976 = w40977 ^ w41015;
	assign w40972 = w40976 ^ w45092;
	assign w40971 = w40995 ^ w40972;
	assign w45983 = w40970 ^ w40971;
	assign w40975 = w41014 ^ w40972;
	assign w41079 = w40974 ^ w40975;
	assign w45986 = ~w41079;
	assign w50935 = w45986 ^ w844;
	assign w50932 = w45983 ^ w841;
	assign w39712 = w39671 ^ w39662;
	assign w39708 = w39712 & w39711;
	assign w39703 = w39708 ^ w39668;
	assign w42135 = w42060 ^ w42150;
	assign w42126 = w42150 & w42135;
	assign w42078 = w42126 ^ w45133;
	assign w42035 = w42126 ^ w42127;
	assign w42082 = w42035 ^ w42036;
	assign w42081 = w42082 ^ w42064;
	assign w42146 = w46159 ^ w42066;
	assign w42142 = w46163 ^ w42146;
	assign w42129 = w42146 & w42142;
	assign w42034 = w42129 ^ w42078;
	assign w42116 = w46163 ^ w42034;
	assign w45061 = w40383 ^ w40389;
	assign w40295 = w40327 ^ w45061;
	assign w40338 = w46143 ^ w40295;
	assign w40333 = w45061 ^ w40318;
	assign w42123 = w42129 ^ w42081;
	assign w42139 = w46164 ^ w42140;
	assign w42132 = w42141 & w42139;
	assign w42083 = w42126 ^ w42132;
	assign w42124 = w42083 ^ w42074;
	assign w42120 = w42124 & w42123;
	assign w42119 = w42120 ^ w42122;
	assign w42121 = w42083 ^ w42075;
	assign w42118 = w42121 & w42119;
	assign w42026 = w42118 ^ w42074;
	assign w42029 = w42118 ^ w42130;
	assign w42025 = w42029 ^ w42065;
	assign w42024 = w46159 ^ w42025;
	assign w42028 = w46157 ^ w42025;
	assign w42115 = w42120 ^ w42080;
	assign w42114 = w42115 & w42116;
	assign w42112 = w42120 ^ w42114;
	assign w42111 = w42122 & w42112;
	assign w42032 = w42114 ^ w42131;
	assign w42027 = w42032 ^ w42128;
	assign w42105 = w42027 ^ w42028;
	assign w42086 = w42105 & w42148;
	assign w42095 = w42105 & w42137;
	assign w42109 = w42111 ^ w42119;
	assign w42033 = w42114 ^ w42078;
	assign w45135 = w42111 ^ w42129;
	assign w42070 = w46163 ^ w45135;
	assign w42110 = w42070 ^ w42033;
	assign w42100 = w42110 & w42139;
	assign w42091 = w42110 & w42141;
	assign w42103 = w45135 ^ w42081;
	assign w42092 = w42103 & w42144;
	assign w42101 = w42103 & w42140;
	assign w42113 = w42114 ^ w42122;
	assign w42090 = w42113 & w42145;
	assign w42099 = w42113 & w46164;
	assign w45138 = w42099 ^ w42101;
	assign w40390 = w40399 & w40397;
	assign w40341 = w40384 ^ w40390;
	assign w40379 = w40341 ^ w40333;
	assign w40382 = w40341 ^ w40332;
	assign w40378 = w40382 & w40381;
	assign w40377 = w40378 ^ w40380;
	assign w40376 = w40379 & w40377;
	assign w40284 = w40376 ^ w40332;
	assign w40287 = w40376 ^ w40388;
	assign w40375 = w40376 ^ w40338;
	assign w40354 = w40375 & w40394;
	assign w40373 = w40378 ^ w40338;
	assign w40372 = w40373 & w40374;
	assign w40370 = w40378 ^ w40372;
	assign w40369 = w40380 & w40370;
	assign w40371 = w40372 ^ w40380;
	assign w40348 = w40371 & w40403;
	assign w40291 = w40372 ^ w40336;
	assign w40290 = w40372 ^ w40389;
	assign w40357 = w40371 & w46148;
	assign w40345 = w40375 & w40401;
	assign w40283 = w40287 ^ w40323;
	assign w40282 = w46143 ^ w40283;
	assign w40367 = w40369 ^ w40377;
	assign w40366 = w40375 & w40367;
	assign w40331 = w40366 ^ w40341;
	assign w40362 = w40331 ^ w40284;
	assign w40347 = w40362 & w40407;
	assign w40289 = w40366 ^ w40390;
	assign w40286 = w46141 ^ w40283;
	assign w45065 = w40369 ^ w40387;
	assign w40361 = w45065 ^ w40339;
	assign w40350 = w40361 & w40402;
	assign w40359 = w40361 & w40398;
	assign w45064 = w40357 ^ w40359;
	assign w40328 = w46147 ^ w45065;
	assign w40368 = w40328 ^ w40291;
	assign w40358 = w40368 & w40397;
	assign w40356 = w40362 & w40392;
	assign w40314 = w40356 ^ w40347;
	assign w40285 = w40290 ^ w40386;
	assign w40365 = w40331 ^ w40333;
	assign w40346 = w40365 & w40400;
	assign w40316 = w40354 ^ w40346;
	assign w40355 = w40365 & w40404;
	assign w40298 = w40354 ^ w40355;
	assign w45063 = w40355 ^ w40356;
	assign w40349 = w40368 & w40399;
	assign w40281 = w40328 ^ w40289;
	assign w40288 = w40318 ^ w40281;
	assign w40364 = w40285 ^ w40288;
	assign w40342 = w40364 & w40405;
	assign w40351 = w40364 & w40396;
	assign w40329 = w40347 ^ w40351;
	assign w40307 = ~w40329;
	assign w40360 = w40281 ^ w40282;
	assign w40352 = w40360 & w40393;
	assign w40337 = w40352 ^ w45063;
	assign w40303 = w40348 ^ w40337;
	assign w40300 = ~w40303;
	assign w40313 = w40352 ^ w40355;
	assign w40310 = ~w40313;
	assign w40343 = w40360 & w40408;
	assign w40306 = w40307 ^ w40345;
	assign w40302 = w40306 ^ w45064;
	assign w40363 = w40285 ^ w40286;
	assign w40353 = w40363 & w40395;
	assign w40297 = w40353 ^ w40337;
	assign w40308 = w40353 ^ w40342;
	assign w40304 = ~w40308;
	assign w40309 = w40352 ^ w40353;
	assign w40344 = w40363 & w40406;
	assign w40305 = w40344 ^ w40302;
	assign w40409 = w40304 ^ w40305;
	assign w46090 = ~w40409;
	assign w51039 = w46090 ^ w756;
	assign w43610 = w40343 ^ w40344;
	assign w40325 = w40349 ^ w43610;
	assign w40326 = w40350 ^ w40325;
	assign w46092 = w40326 ^ w40297;
	assign w40330 = w40358 ^ w40326;
	assign w40299 = w40357 ^ w40330;
	assign w46088 = w40298 ^ w40299;
	assign w40335 = w40359 ^ w40330;
	assign w40410 = w40335 ^ w40309;
	assign w46091 = ~w40410;
	assign w46089 = w45063 ^ w40335;
	assign w51038 = w46089 ^ w755;
	assign w51037 = w46088 ^ w754;
	assign w40312 = w40316 ^ w43610;
	assign w40311 = w40307 ^ w40312;
	assign w40411 = w40310 ^ w40311;
	assign w46086 = ~w40411;
	assign w51035 = w46086 ^ w752;
	assign w51040 = w46091 ^ w757;
	assign w51041 = w46092 ^ w758;
	assign w40315 = w45064 ^ w40312;
	assign w40412 = w40314 ^ w40315;
	assign w46085 = ~w40412;
	assign w51034 = w46085 ^ w751;
	assign w40301 = w40325 ^ w40302;
	assign w46087 = w40300 ^ w40301;
	assign w51036 = w46087 ^ w753;
	assign w39724 = w39654 ^ w39649;
	assign w39716 = w39731 & w39724;
	assign w45033 = w39713 ^ w39716;
	assign w39626 = w39652 ^ w45033;
	assign w39710 = w39626 ^ w39651;
	assign w39666 = w39714 ^ w45033;
	assign w39622 = w39717 ^ w39666;
	assign w39704 = w46139 ^ w39622;
	assign w39707 = w39708 ^ w39710;
	assign w39702 = w39703 & w39704;
	assign w39701 = w39702 ^ w39710;
	assign w39700 = w39708 ^ w39702;
	assign w39699 = w39710 & w39700;
	assign w39697 = w39699 ^ w39707;
	assign w45037 = w39699 ^ w39717;
	assign w39658 = w46139 ^ w45037;
	assign w39678 = w39701 & w39733;
	assign w39620 = w39702 ^ w39719;
	assign w39615 = w39620 ^ w39716;
	assign w39687 = w39701 & w46140;
	assign w39621 = w39702 ^ w39666;
	assign w39698 = w39658 ^ w39621;
	assign w39679 = w39698 & w39729;
	assign w39688 = w39698 & w39727;
	assign w39706 = w39709 & w39707;
	assign w39617 = w39706 ^ w39718;
	assign w39705 = w39706 ^ w39668;
	assign w39696 = w39705 & w39697;
	assign w39619 = w39696 ^ w39720;
	assign w39613 = w39617 ^ w39653;
	assign w39684 = w39705 & w39724;
	assign w39614 = w39706 ^ w39662;
	assign w39675 = w39705 & w39731;
	assign w39612 = w46135 ^ w39613;
	assign w39611 = w39658 ^ w39619;
	assign w39618 = w39648 ^ w39611;
	assign w39694 = w39615 ^ w39618;
	assign w39681 = w39694 & w39726;
	assign w39672 = w39694 & w39735;
	assign w39690 = w39611 ^ w39612;
	assign w39673 = w39690 & w39738;
	assign w39682 = w39690 & w39723;
	assign w39691 = w45037 ^ w39669;
	assign w39680 = w39691 & w39732;
	assign w39689 = w39691 & w39728;
	assign w45036 = w39687 ^ w39689;
	assign w39616 = w46133 ^ w39613;
	assign w39693 = w39615 ^ w39616;
	assign w39674 = w39693 & w39736;
	assign w45034 = w39673 ^ w39674;
	assign w39655 = w39679 ^ w45034;
	assign w39656 = w39680 ^ w39655;
	assign w39660 = w39688 ^ w39656;
	assign w39665 = w39689 ^ w39660;
	assign w39629 = w39687 ^ w39660;
	assign w39683 = w39693 & w39725;
	assign w39639 = w39682 ^ w39683;
	assign w39740 = w39665 ^ w39639;
	assign w46067 = ~w39740;
	assign w51016 = w46067 ^ w797;
	assign w39661 = w39696 ^ w39671;
	assign w39695 = w39661 ^ w39663;
	assign w39685 = w39695 & w39734;
	assign w39692 = w39661 ^ w39614;
	assign w39677 = w39692 & w39737;
	assign w39659 = w39677 ^ w39681;
	assign w39676 = w39695 & w39730;
	assign w39637 = ~w39659;
	assign w39646 = w39684 ^ w39676;
	assign w39643 = w39682 ^ w39685;
	assign w39640 = ~w39643;
	assign w39628 = w39684 ^ w39685;
	assign w46064 = w39628 ^ w39629;
	assign w51013 = w46064 ^ w794;
	assign w39636 = w39637 ^ w39675;
	assign w39632 = w39636 ^ w45036;
	assign w39631 = w39655 ^ w39632;
	assign w39635 = w39674 ^ w39632;
	assign w39686 = w39692 & w39722;
	assign w39644 = w39686 ^ w39677;
	assign w39638 = w39683 ^ w39672;
	assign w39634 = ~w39638;
	assign w39739 = w39634 ^ w39635;
	assign w46066 = ~w39739;
	assign w51015 = w46066 ^ w796;
	assign w39642 = w39646 ^ w45034;
	assign w39641 = w39637 ^ w39642;
	assign w39645 = w45036 ^ w39642;
	assign w39742 = w39644 ^ w39645;
	assign w46061 = ~w39742;
	assign w51010 = w46061 ^ w791;
	assign w39741 = w39640 ^ w39641;
	assign w46062 = ~w39741;
	assign w51011 = w46062 ^ w792;
	assign w45035 = w39685 ^ w39686;
	assign w46065 = w45035 ^ w39665;
	assign w51014 = w46065 ^ w795;
	assign w39667 = w39682 ^ w45035;
	assign w39633 = w39678 ^ w39667;
	assign w39630 = ~w39633;
	assign w46063 = w39630 ^ w39631;
	assign w51012 = w46063 ^ w793;
	assign w39627 = w39683 ^ w39667;
	assign w46068 = w39656 ^ w39627;
	assign w51017 = w46068 ^ w798;
	assign w42117 = w42118 ^ w42080;
	assign w42096 = w42117 & w42136;
	assign w42108 = w42117 & w42109;
	assign w42087 = w42117 & w42143;
	assign w42031 = w42108 ^ w42132;
	assign w42023 = w42070 ^ w42031;
	assign w42030 = w42060 ^ w42023;
	assign w42102 = w42023 ^ w42024;
	assign w42094 = w42102 & w42135;
	assign w42051 = w42094 ^ w42095;
	assign w42106 = w42027 ^ w42030;
	assign w42093 = w42106 & w42138;
	assign w42084 = w42106 & w42147;
	assign w42073 = w42108 ^ w42083;
	assign w42107 = w42073 ^ w42075;
	assign w42088 = w42107 & w42142;
	assign w42104 = w42073 ^ w42026;
	assign w42098 = w42104 & w42134;
	assign w42089 = w42104 & w42149;
	assign w42071 = w42089 ^ w42093;
	assign w42049 = ~w42071;
	assign w42048 = w42049 ^ w42087;
	assign w42044 = w42048 ^ w45138;
	assign w42047 = w42086 ^ w42044;
	assign w42056 = w42098 ^ w42089;
	assign w42097 = w42107 & w42146;
	assign w45137 = w42097 ^ w42098;
	assign w42055 = w42094 ^ w42097;
	assign w42040 = w42096 ^ w42097;
	assign w42079 = w42094 ^ w45137;
	assign w42045 = w42090 ^ w42079;
	assign w42042 = ~w42045;
	assign w42039 = w42095 ^ w42079;
	assign w42085 = w42102 & w42150;
	assign w45134 = w42085 ^ w42086;
	assign w42067 = w42091 ^ w45134;
	assign w42043 = w42067 ^ w42044;
	assign w46007 = w42042 ^ w42043;
	assign w50956 = w46007 ^ w801;
	assign w42068 = w42092 ^ w42067;
	assign w46012 = w42068 ^ w42039;
	assign w42072 = w42100 ^ w42068;
	assign w42041 = w42099 ^ w42072;
	assign w46008 = w42040 ^ w42041;
	assign w50957 = w46008 ^ w802;
	assign w50961 = w46012 ^ w806;
	assign w42050 = w42095 ^ w42084;
	assign w42046 = ~w42050;
	assign w42151 = w42046 ^ w42047;
	assign w46010 = ~w42151;
	assign w50959 = w46010 ^ w804;
	assign w42058 = w42096 ^ w42088;
	assign w42054 = w42058 ^ w45134;
	assign w42057 = w45138 ^ w42054;
	assign w42053 = w42049 ^ w42054;
	assign w42154 = w42056 ^ w42057;
	assign w46005 = ~w42154;
	assign w50954 = w46005 ^ w799;
	assign w42052 = ~w42055;
	assign w42153 = w42052 ^ w42053;
	assign w46006 = ~w42153;
	assign w50955 = w46006 ^ w800;
	assign w3460 = w3471 & w3512;
	assign w3436 = w3460 ^ w3435;
	assign w46100 = w3436 ^ w3407;
	assign w51049 = w46100 ^ w766;
	assign w3440 = w3468 ^ w3436;
	assign w3409 = w3467 ^ w3440;
	assign w46096 = w3408 ^ w3409;
	assign w51045 = w46096 ^ w762;
	assign w3445 = w3469 ^ w3440;
	assign w46097 = w43680 ^ w3445;
	assign w51046 = w46097 ^ w763;
	assign w3520 = w3445 ^ w3419;
	assign w46099 = ~w3520;
	assign w51048 = w46099 ^ w765;
	assign w43649 = w2823 ^ w2826;
	assign w2736 = w2762 ^ w43649;
	assign w2820 = w2736 ^ w2761;
	assign w2817 = w2818 ^ w2820;
	assign w2816 = w2819 & w2817;
	assign w2815 = w2816 ^ w2778;
	assign w2785 = w2815 & w2841;
	assign w2794 = w2815 & w2834;
	assign w2727 = w2816 ^ w2828;
	assign w2723 = w2727 ^ w2763;
	assign w2726 = w46181 ^ w2723;
	assign w2722 = w46183 ^ w2723;
	assign w2724 = w2816 ^ w2772;
	assign w2776 = w2824 ^ w43649;
	assign w2732 = w2827 ^ w2776;
	assign w2814 = w46187 ^ w2732;
	assign w2812 = w2813 & w2814;
	assign w2810 = w2818 ^ w2812;
	assign w2809 = w2820 & w2810;
	assign w2811 = w2812 ^ w2820;
	assign w2788 = w2811 & w2843;
	assign w2797 = w2811 & w46188;
	assign w2807 = w2809 ^ w2817;
	assign w2806 = w2815 & w2807;
	assign w2729 = w2806 ^ w2830;
	assign w2731 = w2812 ^ w2776;
	assign w43652 = w2809 ^ w2827;
	assign w2801 = w43652 ^ w2779;
	assign w2790 = w2801 & w2842;
	assign w2768 = w46187 ^ w43652;
	assign w2721 = w2768 ^ w2729;
	assign w2800 = w2721 ^ w2722;
	assign w2792 = w2800 & w2833;
	assign w2783 = w2800 & w2848;
	assign w2808 = w2768 ^ w2731;
	assign w2789 = w2808 & w2839;
	assign w2798 = w2808 & w2837;
	assign w2771 = w2806 ^ w2781;
	assign w2805 = w2771 ^ w2773;
	assign w2795 = w2805 & w2844;
	assign w2738 = w2794 ^ w2795;
	assign w2753 = w2792 ^ w2795;
	assign w2786 = w2805 & w2840;
	assign w2750 = ~w2753;
	assign w2730 = w2812 ^ w2829;
	assign w2725 = w2730 ^ w2826;
	assign w2803 = w2725 ^ w2726;
	assign w2793 = w2803 & w2835;
	assign w2749 = w2792 ^ w2793;
	assign w2784 = w2803 & w2846;
	assign w43514 = w2783 ^ w2784;
	assign w2765 = w2789 ^ w43514;
	assign w2756 = w2794 ^ w2786;
	assign w2752 = w2756 ^ w43514;
	assign w2728 = w2758 ^ w2721;
	assign w2804 = w2725 ^ w2728;
	assign w2782 = w2804 & w2845;
	assign w2748 = w2793 ^ w2782;
	assign w2791 = w2804 & w2836;
	assign w2744 = ~w2748;
	assign w2799 = w2801 & w2838;
	assign w43651 = w2797 ^ w2799;
	assign w2755 = w43651 ^ w2752;
	assign w2766 = w2790 ^ w2765;
	assign w2770 = w2798 ^ w2766;
	assign w2775 = w2799 ^ w2770;
	assign w2739 = w2797 ^ w2770;
	assign w2850 = w2775 ^ w2749;
	assign w46083 = ~w2850;
	assign w46080 = w2738 ^ w2739;
	assign w51029 = w46080 ^ w746;
	assign w51032 = w46083 ^ w749;
	assign w2802 = w2771 ^ w2724;
	assign w2796 = w2802 & w2832;
	assign w2787 = w2802 & w2847;
	assign w2769 = w2787 ^ w2791;
	assign w2754 = w2796 ^ w2787;
	assign w2852 = w2754 ^ w2755;
	assign w2747 = ~w2769;
	assign w2746 = w2747 ^ w2785;
	assign w2742 = w2746 ^ w43651;
	assign w2741 = w2765 ^ w2742;
	assign w2751 = w2747 ^ w2752;
	assign w2851 = w2750 ^ w2751;
	assign w46078 = ~w2851;
	assign w2745 = w2784 ^ w2742;
	assign w2849 = w2744 ^ w2745;
	assign w51027 = w46078 ^ w744;
	assign w46082 = ~w2849;
	assign w51031 = w46082 ^ w748;
	assign w46077 = ~w2852;
	assign w51026 = w46077 ^ w743;
	assign w43650 = w2795 ^ w2796;
	assign w2777 = w2792 ^ w43650;
	assign w2743 = w2788 ^ w2777;
	assign w2740 = ~w2743;
	assign w46079 = w2740 ^ w2741;
	assign w51028 = w46079 ^ w745;
	assign w2737 = w2793 ^ w2777;
	assign w46084 = w2766 ^ w2737;
	assign w51033 = w46084 ^ w750;
	assign w46081 = w43650 ^ w2775;
	assign w51030 = w46081 ^ w747;
	assign w42077 = w42101 ^ w42072;
	assign w42152 = w42077 ^ w42051;
	assign w46009 = w45137 ^ w42077;
	assign w50958 = w46009 ^ w803;
	assign w46011 = ~w42152;
	assign w50960 = w46011 ^ w805;
	assign w42190 = w42232 ^ w42223;
	assign w42288 = w42190 ^ w42191;
	assign w46053 = ~w42288;
	assign w51002 = w46053 ^ w783;
	assign w2912 = w46167 ^ w2869;
	assign w50835 = w10408 ^ w10409;
	assign w46114 = w50835 ^ w625;
	assign w3270 = w46113 ^ w46114;
	assign w3295 = w46114 ^ w3293;
	assign w3368 = w46111 ^ w3295;
	assign w3370 = w3300 ^ w3295;
	assign w3364 = w3383 & w3368;
	assign w3298 = w3364 ^ w3294;
	assign w3310 = w46115 ^ w46114;
	assign w3378 = w3382 ^ w3310;
	assign w3367 = w3374 & w3378;
	assign w3384 = w46114 ^ w46112;
	assign w3369 = w3294 ^ w3384;
	assign w3360 = w3384 & w3369;
	assign w3362 = w3377 & w3370;
	assign w3375 = w3310 ^ w3377;
	assign w3366 = w3375 & w3373;
	assign w3317 = w3360 ^ w3366;
	assign w3299 = w3367 ^ w3296;
	assign w3381 = w46109 ^ w46114;
	assign w3359 = w3381 & w3372;
	assign w43670 = w3359 ^ w3365;
	assign w3309 = w43670 ^ w3294;
	assign w3355 = w3317 ^ w3309;
	assign w43671 = w3359 ^ w3362;
	assign w3272 = w3298 ^ w43671;
	assign w3312 = w3360 ^ w43671;
	assign w3268 = w3363 ^ w3312;
	assign w3350 = w46115 ^ w3268;
	assign w3371 = w46110 ^ w3295;
	assign w3361 = w3382 & w3371;
	assign w3269 = w3360 ^ w3361;
	assign w3316 = w3269 ^ w3270;
	assign w3315 = w3316 ^ w3298;
	assign w3357 = w3363 ^ w3315;
	assign w3297 = w3361 ^ w3295;
	assign w3303 = w3299 ^ w3297;
	assign w3356 = w3272 ^ w3297;
	assign w3308 = w46109 ^ w3303;
	assign w3358 = w3317 ^ w3308;
	assign w3271 = w3303 ^ w43670;
	assign w3314 = w46111 ^ w3271;
	assign w3354 = w3358 & w3357;
	assign w3353 = w3354 ^ w3356;
	assign w3349 = w3354 ^ w3314;
	assign w3348 = w3349 & w3350;
	assign w3267 = w3348 ^ w3312;
	assign w3266 = w3348 ^ w3365;
	assign w3261 = w3266 ^ w3362;
	assign w3347 = w3348 ^ w3356;
	assign w3324 = w3347 & w3379;
	assign w3333 = w3347 & w46116;
	assign w3346 = w3354 ^ w3348;
	assign w3352 = w3355 & w3353;
	assign w3260 = w3352 ^ w3308;
	assign w3351 = w3352 ^ w3314;
	assign w3321 = w3351 & w3377;
	assign w3330 = w3351 & w3370;
	assign w3263 = w3352 ^ w3364;
	assign w3259 = w3263 ^ w3299;
	assign w3262 = w46109 ^ w3259;
	assign w3258 = w46111 ^ w3259;
	assign w3339 = w3261 ^ w3262;
	assign w3329 = w3339 & w3371;
	assign w3320 = w3339 & w3382;
	assign w3345 = w3356 & w3346;
	assign w3343 = w3345 ^ w3353;
	assign w3342 = w3351 & w3343;
	assign w3307 = w3342 ^ w3317;
	assign w3338 = w3307 ^ w3260;
	assign w3332 = w3338 & w3368;
	assign w3323 = w3338 & w3383;
	assign w3290 = w3332 ^ w3323;
	assign w3265 = w3342 ^ w3366;
	assign w3341 = w3307 ^ w3309;
	assign w3322 = w3341 & w3376;
	assign w3292 = w3330 ^ w3322;
	assign w3331 = w3341 & w3380;
	assign w43673 = w3331 ^ w3332;
	assign w3274 = w3330 ^ w3331;
	assign w43675 = w3345 ^ w3363;
	assign w3337 = w43675 ^ w3315;
	assign w3335 = w3337 & w3374;
	assign w43674 = w3333 ^ w3335;
	assign w3326 = w3337 & w3378;
	assign w3304 = w46115 ^ w43675;
	assign w3257 = w3304 ^ w3265;
	assign w3264 = w3294 ^ w3257;
	assign w3340 = w3261 ^ w3264;
	assign w3318 = w3340 & w3381;
	assign w3327 = w3340 & w3372;
	assign w3305 = w3323 ^ w3327;
	assign w3283 = ~w3305;
	assign w3282 = w3283 ^ w3321;
	assign w3284 = w3329 ^ w3318;
	assign w3344 = w3304 ^ w3267;
	assign w3325 = w3344 & w3375;
	assign w3334 = w3344 & w3373;
	assign w3278 = w3282 ^ w43674;
	assign w3281 = w3320 ^ w3278;
	assign w3336 = w3257 ^ w3258;
	assign w3319 = w3336 & w3384;
	assign w43672 = w3319 ^ w3320;
	assign w3301 = w3325 ^ w43672;
	assign w3302 = w3326 ^ w3301;
	assign w3306 = w3334 ^ w3302;
	assign w3328 = w3336 & w3369;
	assign w3289 = w3328 ^ w3331;
	assign w3286 = ~w3289;
	assign w3313 = w3328 ^ w43673;
	assign w3279 = w3324 ^ w3313;
	assign w3285 = w3328 ^ w3329;
	assign w3288 = w3292 ^ w43672;
	assign w3291 = w43674 ^ w3288;
	assign w3388 = w3290 ^ w3291;
	assign w3287 = w3283 ^ w3288;
	assign w3387 = w3286 ^ w3287;
	assign w45989 = ~w3388;
	assign w50938 = w45989 ^ w847;
	assign w45990 = ~w3387;
	assign w50939 = w45990 ^ w848;
	assign w3311 = w3335 ^ w3306;
	assign w45993 = w43673 ^ w3311;
	assign w3386 = w3311 ^ w3285;
	assign w45995 = ~w3386;
	assign w50944 = w45995 ^ w853;
	assign w3273 = w3329 ^ w3313;
	assign w3275 = w3333 ^ w3306;
	assign w45992 = w3274 ^ w3275;
	assign w50941 = w45992 ^ w850;
	assign w45996 = w3302 ^ w3273;
	assign w50945 = w45996 ^ w854;
	assign w3276 = ~w3279;
	assign w50942 = w45993 ^ w851;
	assign w3277 = w3301 ^ w3278;
	assign w45991 = w3276 ^ w3277;
	assign w50940 = w45991 ^ w849;
	assign w3280 = ~w3284;
	assign w3385 = w3280 ^ w3281;
	assign w45994 = ~w3385;
	assign w50943 = w45994 ^ w852;
	assign w2256 = w2264 & w2297;
	assign w2213 = w2256 ^ w2257;
	assign w2314 = w2239 ^ w2213;
	assign w2241 = w2256 ^ w43629;
	assign w2201 = w2257 ^ w2241;
	assign w2207 = w2252 ^ w2241;
	assign w46052 = w2230 ^ w2201;
	assign w51001 = w46052 ^ w782;
	assign w2217 = w2256 ^ w2259;
	assign w46051 = ~w2314;
	assign w51000 = w46051 ^ w781;
	assign w2214 = ~w2217;
	assign w2315 = w2214 ^ w2215;
	assign w46046 = ~w2315;
	assign w50995 = w46046 ^ w776;
	assign w2204 = ~w2207;
	assign w46047 = w2204 ^ w2205;
	assign w50996 = w46047 ^ w777;
	assign w2914 = w2867 ^ w2868;
	assign w2913 = w2914 ^ w2896;
	assign w2955 = w2961 ^ w2913;
	assign w2952 = w2956 & w2955;
	assign w2951 = w2952 ^ w2954;
	assign w2947 = w2952 ^ w2912;
	assign w2946 = w2947 & w2948;
	assign w2945 = w2946 ^ w2954;
	assign w2922 = w2945 & w2977;
	assign w2944 = w2952 ^ w2946;
	assign w2943 = w2954 & w2944;
	assign w43658 = w2943 ^ w2961;
	assign w2935 = w43658 ^ w2913;
	assign w2924 = w2935 & w2976;
	assign w2902 = w46171 ^ w43658;
	assign w2950 = w2953 & w2951;
	assign w2861 = w2950 ^ w2962;
	assign w2949 = w2950 ^ w2912;
	assign w2919 = w2949 & w2975;
	assign w2933 = w2935 & w2972;
	assign w2858 = w2950 ^ w2906;
	assign w2928 = w2949 & w2968;
	assign w2941 = w2943 ^ w2951;
	assign w2940 = w2949 & w2941;
	assign w2863 = w2940 ^ w2964;
	assign w2905 = w2940 ^ w2915;
	assign w2939 = w2905 ^ w2907;
	assign w2929 = w2939 & w2978;
	assign w2872 = w2928 ^ w2929;
	assign w2936 = w2905 ^ w2858;
	assign w2921 = w2936 & w2981;
	assign w2930 = w2936 & w2966;
	assign w43656 = w2929 ^ w2930;
	assign w2888 = w2930 ^ w2921;
	assign w2931 = w2945 & w46172;
	assign w43657 = w2931 ^ w2933;
	assign w2920 = w2939 & w2974;
	assign w2890 = w2928 ^ w2920;
	assign w2865 = w2946 ^ w2910;
	assign w2942 = w2902 ^ w2865;
	assign w2923 = w2942 & w2973;
	assign w2932 = w2942 & w2971;
	assign w2857 = w2861 ^ w2897;
	assign w2860 = w46165 ^ w2857;
	assign w2856 = w46167 ^ w2857;
	assign w2864 = w2946 ^ w2963;
	assign w2859 = w2864 ^ w2960;
	assign w2937 = w2859 ^ w2860;
	assign w2918 = w2937 & w2980;
	assign w2927 = w2937 & w2969;
	assign w2855 = w2902 ^ w2863;
	assign w2862 = w2892 ^ w2855;
	assign w2938 = w2859 ^ w2862;
	assign w2916 = w2938 & w2979;
	assign w2882 = w2927 ^ w2916;
	assign w2878 = ~w2882;
	assign w2925 = w2938 & w2970;
	assign w2903 = w2921 ^ w2925;
	assign w2881 = ~w2903;
	assign w2880 = w2881 ^ w2919;
	assign w2934 = w2855 ^ w2856;
	assign w2917 = w2934 & w2982;
	assign w2926 = w2934 & w2967;
	assign w2887 = w2926 ^ w2929;
	assign w2884 = ~w2887;
	assign w2911 = w2926 ^ w43656;
	assign w2877 = w2922 ^ w2911;
	assign w2883 = w2926 ^ w2927;
	assign w2871 = w2927 ^ w2911;
	assign w2874 = ~w2877;
	assign w43655 = w2917 ^ w2918;
	assign w2886 = w2890 ^ w43655;
	assign w2885 = w2881 ^ w2886;
	assign w2985 = w2884 ^ w2885;
	assign w2899 = w2923 ^ w43655;
	assign w2900 = w2924 ^ w2899;
	assign w46036 = w2900 ^ w2871;
	assign w50985 = w46036 ^ w830;
	assign w2904 = w2932 ^ w2900;
	assign w2873 = w2931 ^ w2904;
	assign w2909 = w2933 ^ w2904;
	assign w2984 = w2909 ^ w2883;
	assign w46035 = ~w2984;
	assign w50984 = w46035 ^ w829;
	assign w2889 = w43657 ^ w2886;
	assign w2986 = w2888 ^ w2889;
	assign w46029 = ~w2986;
	assign w50978 = w46029 ^ w823;
	assign w46033 = w43656 ^ w2909;
	assign w50982 = w46033 ^ w827;
	assign w46032 = w2872 ^ w2873;
	assign w50981 = w46032 ^ w826;
	assign w46030 = ~w2985;
	assign w50979 = w46030 ^ w824;
	assign w2876 = w2880 ^ w43657;
	assign w2879 = w2918 ^ w2876;
	assign w2983 = w2878 ^ w2879;
	assign w46034 = ~w2983;
	assign w50983 = w46034 ^ w828;
	assign w2875 = w2899 ^ w2876;
	assign w46031 = w2874 ^ w2875;
	assign w50980 = w46031 ^ w825;

endmodule
