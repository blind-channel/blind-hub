module sha256(
    input wire [511:0] data,
    input wire [255:0] state,
    output wire [255:0] next_state,
);
    raw_sha256 sha(
        .w0(data[0]),
        .w1(data[1]),
        .w2(data[2]),
        .w3(data[3]),
        .w4(data[4]),
        .w5(data[5]),
        .w6(data[6]),
        .w7(data[7]),
        .w8(data[8]),
        .w9(data[9]),
        .w10(data[10]),
        .w11(data[11]),
        .w12(data[12]),
        .w13(data[13]),
        .w14(data[14]),
        .w15(data[15]),
        .w16(data[16]),
        .w17(data[17]),
        .w18(data[18]),
        .w19(data[19]),
        .w20(data[20]),
        .w21(data[21]),
        .w22(data[22]),
        .w23(data[23]),
        .w24(data[24]),
        .w25(data[25]),
        .w26(data[26]),
        .w27(data[27]),
        .w28(data[28]),
        .w29(data[29]),
        .w30(data[30]),
        .w31(data[31]),
        .w32(data[32]),
        .w33(data[33]),
        .w34(data[34]),
        .w35(data[35]),
        .w36(data[36]),
        .w37(data[37]),
        .w38(data[38]),
        .w39(data[39]),
        .w40(data[40]),
        .w41(data[41]),
        .w42(data[42]),
        .w43(data[43]),
        .w44(data[44]),
        .w45(data[45]),
        .w46(data[46]),
        .w47(data[47]),
        .w48(data[48]),
        .w49(data[49]),
        .w50(data[50]),
        .w51(data[51]),
        .w52(data[52]),
        .w53(data[53]),
        .w54(data[54]),
        .w55(data[55]),
        .w56(data[56]),
        .w57(data[57]),
        .w58(data[58]),
        .w59(data[59]),
        .w60(data[60]),
        .w61(data[61]),
        .w62(data[62]),
        .w63(data[63]),
        .w64(data[64]),
        .w65(data[65]),
        .w66(data[66]),
        .w67(data[67]),
        .w68(data[68]),
        .w69(data[69]),
        .w70(data[70]),
        .w71(data[71]),
        .w72(data[72]),
        .w73(data[73]),
        .w74(data[74]),
        .w75(data[75]),
        .w76(data[76]),
        .w77(data[77]),
        .w78(data[78]),
        .w79(data[79]),
        .w80(data[80]),
        .w81(data[81]),
        .w82(data[82]),
        .w83(data[83]),
        .w84(data[84]),
        .w85(data[85]),
        .w86(data[86]),
        .w87(data[87]),
        .w88(data[88]),
        .w89(data[89]),
        .w90(data[90]),
        .w91(data[91]),
        .w92(data[92]),
        .w93(data[93]),
        .w94(data[94]),
        .w95(data[95]),
        .w96(data[96]),
        .w97(data[97]),
        .w98(data[98]),
        .w99(data[99]),
        .w100(data[100]),
        .w101(data[101]),
        .w102(data[102]),
        .w103(data[103]),
        .w104(data[104]),
        .w105(data[105]),
        .w106(data[106]),
        .w107(data[107]),
        .w108(data[108]),
        .w109(data[109]),
        .w110(data[110]),
        .w111(data[111]),
        .w112(data[112]),
        .w113(data[113]),
        .w114(data[114]),
        .w115(data[115]),
        .w116(data[116]),
        .w117(data[117]),
        .w118(data[118]),
        .w119(data[119]),
        .w120(data[120]),
        .w121(data[121]),
        .w122(data[122]),
        .w123(data[123]),
        .w124(data[124]),
        .w125(data[125]),
        .w126(data[126]),
        .w127(data[127]),
        .w128(data[128]),
        .w129(data[129]),
        .w130(data[130]),
        .w131(data[131]),
        .w132(data[132]),
        .w133(data[133]),
        .w134(data[134]),
        .w135(data[135]),
        .w136(data[136]),
        .w137(data[137]),
        .w138(data[138]),
        .w139(data[139]),
        .w140(data[140]),
        .w141(data[141]),
        .w142(data[142]),
        .w143(data[143]),
        .w144(data[144]),
        .w145(data[145]),
        .w146(data[146]),
        .w147(data[147]),
        .w148(data[148]),
        .w149(data[149]),
        .w150(data[150]),
        .w151(data[151]),
        .w152(data[152]),
        .w153(data[153]),
        .w154(data[154]),
        .w155(data[155]),
        .w156(data[156]),
        .w157(data[157]),
        .w158(data[158]),
        .w159(data[159]),
        .w160(data[160]),
        .w161(data[161]),
        .w162(data[162]),
        .w163(data[163]),
        .w164(data[164]),
        .w165(data[165]),
        .w166(data[166]),
        .w167(data[167]),
        .w168(data[168]),
        .w169(data[169]),
        .w170(data[170]),
        .w171(data[171]),
        .w172(data[172]),
        .w173(data[173]),
        .w174(data[174]),
        .w175(data[175]),
        .w176(data[176]),
        .w177(data[177]),
        .w178(data[178]),
        .w179(data[179]),
        .w180(data[180]),
        .w181(data[181]),
        .w182(data[182]),
        .w183(data[183]),
        .w184(data[184]),
        .w185(data[185]),
        .w186(data[186]),
        .w187(data[187]),
        .w188(data[188]),
        .w189(data[189]),
        .w190(data[190]),
        .w191(data[191]),
        .w192(data[192]),
        .w193(data[193]),
        .w194(data[194]),
        .w195(data[195]),
        .w196(data[196]),
        .w197(data[197]),
        .w198(data[198]),
        .w199(data[199]),
        .w200(data[200]),
        .w201(data[201]),
        .w202(data[202]),
        .w203(data[203]),
        .w204(data[204]),
        .w205(data[205]),
        .w206(data[206]),
        .w207(data[207]),
        .w208(data[208]),
        .w209(data[209]),
        .w210(data[210]),
        .w211(data[211]),
        .w212(data[212]),
        .w213(data[213]),
        .w214(data[214]),
        .w215(data[215]),
        .w216(data[216]),
        .w217(data[217]),
        .w218(data[218]),
        .w219(data[219]),
        .w220(data[220]),
        .w221(data[221]),
        .w222(data[222]),
        .w223(data[223]),
        .w224(data[224]),
        .w225(data[225]),
        .w226(data[226]),
        .w227(data[227]),
        .w228(data[228]),
        .w229(data[229]),
        .w230(data[230]),
        .w231(data[231]),
        .w232(data[232]),
        .w233(data[233]),
        .w234(data[234]),
        .w235(data[235]),
        .w236(data[236]),
        .w237(data[237]),
        .w238(data[238]),
        .w239(data[239]),
        .w240(data[240]),
        .w241(data[241]),
        .w242(data[242]),
        .w243(data[243]),
        .w244(data[244]),
        .w245(data[245]),
        .w246(data[246]),
        .w247(data[247]),
        .w248(data[248]),
        .w249(data[249]),
        .w250(data[250]),
        .w251(data[251]),
        .w252(data[252]),
        .w253(data[253]),
        .w254(data[254]),
        .w255(data[255]),
        .w256(data[256]),
        .w257(data[257]),
        .w258(data[258]),
        .w259(data[259]),
        .w260(data[260]),
        .w261(data[261]),
        .w262(data[262]),
        .w263(data[263]),
        .w264(data[264]),
        .w265(data[265]),
        .w266(data[266]),
        .w267(data[267]),
        .w268(data[268]),
        .w269(data[269]),
        .w270(data[270]),
        .w271(data[271]),
        .w272(data[272]),
        .w273(data[273]),
        .w274(data[274]),
        .w275(data[275]),
        .w276(data[276]),
        .w277(data[277]),
        .w278(data[278]),
        .w279(data[279]),
        .w280(data[280]),
        .w281(data[281]),
        .w282(data[282]),
        .w283(data[283]),
        .w284(data[284]),
        .w285(data[285]),
        .w286(data[286]),
        .w287(data[287]),
        .w288(data[288]),
        .w289(data[289]),
        .w290(data[290]),
        .w291(data[291]),
        .w292(data[292]),
        .w293(data[293]),
        .w294(data[294]),
        .w295(data[295]),
        .w296(data[296]),
        .w297(data[297]),
        .w298(data[298]),
        .w299(data[299]),
        .w300(data[300]),
        .w301(data[301]),
        .w302(data[302]),
        .w303(data[303]),
        .w304(data[304]),
        .w305(data[305]),
        .w306(data[306]),
        .w307(data[307]),
        .w308(data[308]),
        .w309(data[309]),
        .w310(data[310]),
        .w311(data[311]),
        .w312(data[312]),
        .w313(data[313]),
        .w314(data[314]),
        .w315(data[315]),
        .w316(data[316]),
        .w317(data[317]),
        .w318(data[318]),
        .w319(data[319]),
        .w320(data[320]),
        .w321(data[321]),
        .w322(data[322]),
        .w323(data[323]),
        .w324(data[324]),
        .w325(data[325]),
        .w326(data[326]),
        .w327(data[327]),
        .w328(data[328]),
        .w329(data[329]),
        .w330(data[330]),
        .w331(data[331]),
        .w332(data[332]),
        .w333(data[333]),
        .w334(data[334]),
        .w335(data[335]),
        .w336(data[336]),
        .w337(data[337]),
        .w338(data[338]),
        .w339(data[339]),
        .w340(data[340]),
        .w341(data[341]),
        .w342(data[342]),
        .w343(data[343]),
        .w344(data[344]),
        .w345(data[345]),
        .w346(data[346]),
        .w347(data[347]),
        .w348(data[348]),
        .w349(data[349]),
        .w350(data[350]),
        .w351(data[351]),
        .w352(data[352]),
        .w353(data[353]),
        .w354(data[354]),
        .w355(data[355]),
        .w356(data[356]),
        .w357(data[357]),
        .w358(data[358]),
        .w359(data[359]),
        .w360(data[360]),
        .w361(data[361]),
        .w362(data[362]),
        .w363(data[363]),
        .w364(data[364]),
        .w365(data[365]),
        .w366(data[366]),
        .w367(data[367]),
        .w368(data[368]),
        .w369(data[369]),
        .w370(data[370]),
        .w371(data[371]),
        .w372(data[372]),
        .w373(data[373]),
        .w374(data[374]),
        .w375(data[375]),
        .w376(data[376]),
        .w377(data[377]),
        .w378(data[378]),
        .w379(data[379]),
        .w380(data[380]),
        .w381(data[381]),
        .w382(data[382]),
        .w383(data[383]),
        .w384(data[384]),
        .w385(data[385]),
        .w386(data[386]),
        .w387(data[387]),
        .w388(data[388]),
        .w389(data[389]),
        .w390(data[390]),
        .w391(data[391]),
        .w392(data[392]),
        .w393(data[393]),
        .w394(data[394]),
        .w395(data[395]),
        .w396(data[396]),
        .w397(data[397]),
        .w398(data[398]),
        .w399(data[399]),
        .w400(data[400]),
        .w401(data[401]),
        .w402(data[402]),
        .w403(data[403]),
        .w404(data[404]),
        .w405(data[405]),
        .w406(data[406]),
        .w407(data[407]),
        .w408(data[408]),
        .w409(data[409]),
        .w410(data[410]),
        .w411(data[411]),
        .w412(data[412]),
        .w413(data[413]),
        .w414(data[414]),
        .w415(data[415]),
        .w416(data[416]),
        .w417(data[417]),
        .w418(data[418]),
        .w419(data[419]),
        .w420(data[420]),
        .w421(data[421]),
        .w422(data[422]),
        .w423(data[423]),
        .w424(data[424]),
        .w425(data[425]),
        .w426(data[426]),
        .w427(data[427]),
        .w428(data[428]),
        .w429(data[429]),
        .w430(data[430]),
        .w431(data[431]),
        .w432(data[432]),
        .w433(data[433]),
        .w434(data[434]),
        .w435(data[435]),
        .w436(data[436]),
        .w437(data[437]),
        .w438(data[438]),
        .w439(data[439]),
        .w440(data[440]),
        .w441(data[441]),
        .w442(data[442]),
        .w443(data[443]),
        .w444(data[444]),
        .w445(data[445]),
        .w446(data[446]),
        .w447(data[447]),
        .w448(data[448]),
        .w449(data[449]),
        .w450(data[450]),
        .w451(data[451]),
        .w452(data[452]),
        .w453(data[453]),
        .w454(data[454]),
        .w455(data[455]),
        .w456(data[456]),
        .w457(data[457]),
        .w458(data[458]),
        .w459(data[459]),
        .w460(data[460]),
        .w461(data[461]),
        .w462(data[462]),
        .w463(data[463]),
        .w464(data[464]),
        .w465(data[465]),
        .w466(data[466]),
        .w467(data[467]),
        .w468(data[468]),
        .w469(data[469]),
        .w470(data[470]),
        .w471(data[471]),
        .w472(data[472]),
        .w473(data[473]),
        .w474(data[474]),
        .w475(data[475]),
        .w476(data[476]),
        .w477(data[477]),
        .w478(data[478]),
        .w479(data[479]),
        .w480(data[480]),
        .w481(data[481]),
        .w482(data[482]),
        .w483(data[483]),
        .w484(data[484]),
        .w485(data[485]),
        .w486(data[486]),
        .w487(data[487]),
        .w488(data[488]),
        .w489(data[489]),
        .w490(data[490]),
        .w491(data[491]),
        .w492(data[492]),
        .w493(data[493]),
        .w494(data[494]),
        .w495(data[495]),
        .w496(data[496]),
        .w497(data[497]),
        .w498(data[498]),
        .w499(data[499]),
        .w500(data[500]),
        .w501(data[501]),
        .w502(data[502]),
        .w503(data[503]),
        .w504(data[504]),
        .w505(data[505]),
        .w506(data[506]),
        .w507(data[507]),
        .w508(data[508]),
        .w509(data[509]),
        .w510(data[510]),
        .w511(data[511]),
        .w512(state[0]),
        .w513(state[1]),
        .w514(state[2]),
        .w515(state[3]),
        .w516(state[4]),
        .w517(state[5]),
        .w518(state[6]),
        .w519(state[7]),
        .w520(state[8]),
        .w521(state[9]),
        .w522(state[10]),
        .w523(state[11]),
        .w524(state[12]),
        .w525(state[13]),
        .w526(state[14]),
        .w527(state[15]),
        .w528(state[16]),
        .w529(state[17]),
        .w530(state[18]),
        .w531(state[19]),
        .w532(state[20]),
        .w533(state[21]),
        .w534(state[22]),
        .w535(state[23]),
        .w536(state[24]),
        .w537(state[25]),
        .w538(state[26]),
        .w539(state[27]),
        .w540(state[28]),
        .w541(state[29]),
        .w542(state[30]),
        .w543(state[31]),
        .w544(state[32]),
        .w545(state[33]),
        .w546(state[34]),
        .w547(state[35]),
        .w548(state[36]),
        .w549(state[37]),
        .w550(state[38]),
        .w551(state[39]),
        .w552(state[40]),
        .w553(state[41]),
        .w554(state[42]),
        .w555(state[43]),
        .w556(state[44]),
        .w557(state[45]),
        .w558(state[46]),
        .w559(state[47]),
        .w560(state[48]),
        .w561(state[49]),
        .w562(state[50]),
        .w563(state[51]),
        .w564(state[52]),
        .w565(state[53]),
        .w566(state[54]),
        .w567(state[55]),
        .w568(state[56]),
        .w569(state[57]),
        .w570(state[58]),
        .w571(state[59]),
        .w572(state[60]),
        .w573(state[61]),
        .w574(state[62]),
        .w575(state[63]),
        .w576(state[64]),
        .w577(state[65]),
        .w578(state[66]),
        .w579(state[67]),
        .w580(state[68]),
        .w581(state[69]),
        .w582(state[70]),
        .w583(state[71]),
        .w584(state[72]),
        .w585(state[73]),
        .w586(state[74]),
        .w587(state[75]),
        .w588(state[76]),
        .w589(state[77]),
        .w590(state[78]),
        .w591(state[79]),
        .w592(state[80]),
        .w593(state[81]),
        .w594(state[82]),
        .w595(state[83]),
        .w596(state[84]),
        .w597(state[85]),
        .w598(state[86]),
        .w599(state[87]),
        .w600(state[88]),
        .w601(state[89]),
        .w602(state[90]),
        .w603(state[91]),
        .w604(state[92]),
        .w605(state[93]),
        .w606(state[94]),
        .w607(state[95]),
        .w608(state[96]),
        .w609(state[97]),
        .w610(state[98]),
        .w611(state[99]),
        .w612(state[100]),
        .w613(state[101]),
        .w614(state[102]),
        .w615(state[103]),
        .w616(state[104]),
        .w617(state[105]),
        .w618(state[106]),
        .w619(state[107]),
        .w620(state[108]),
        .w621(state[109]),
        .w622(state[110]),
        .w623(state[111]),
        .w624(state[112]),
        .w625(state[113]),
        .w626(state[114]),
        .w627(state[115]),
        .w628(state[116]),
        .w629(state[117]),
        .w630(state[118]),
        .w631(state[119]),
        .w632(state[120]),
        .w633(state[121]),
        .w634(state[122]),
        .w635(state[123]),
        .w636(state[124]),
        .w637(state[125]),
        .w638(state[126]),
        .w639(state[127]),
        .w640(state[128]),
        .w641(state[129]),
        .w642(state[130]),
        .w643(state[131]),
        .w644(state[132]),
        .w645(state[133]),
        .w646(state[134]),
        .w647(state[135]),
        .w648(state[136]),
        .w649(state[137]),
        .w650(state[138]),
        .w651(state[139]),
        .w652(state[140]),
        .w653(state[141]),
        .w654(state[142]),
        .w655(state[143]),
        .w656(state[144]),
        .w657(state[145]),
        .w658(state[146]),
        .w659(state[147]),
        .w660(state[148]),
        .w661(state[149]),
        .w662(state[150]),
        .w663(state[151]),
        .w664(state[152]),
        .w665(state[153]),
        .w666(state[154]),
        .w667(state[155]),
        .w668(state[156]),
        .w669(state[157]),
        .w670(state[158]),
        .w671(state[159]),
        .w672(state[160]),
        .w673(state[161]),
        .w674(state[162]),
        .w675(state[163]),
        .w676(state[164]),
        .w677(state[165]),
        .w678(state[166]),
        .w679(state[167]),
        .w680(state[168]),
        .w681(state[169]),
        .w682(state[170]),
        .w683(state[171]),
        .w684(state[172]),
        .w685(state[173]),
        .w686(state[174]),
        .w687(state[175]),
        .w688(state[176]),
        .w689(state[177]),
        .w690(state[178]),
        .w691(state[179]),
        .w692(state[180]),
        .w693(state[181]),
        .w694(state[182]),
        .w695(state[183]),
        .w696(state[184]),
        .w697(state[185]),
        .w698(state[186]),
        .w699(state[187]),
        .w700(state[188]),
        .w701(state[189]),
        .w702(state[190]),
        .w703(state[191]),
        .w704(state[192]),
        .w705(state[193]),
        .w706(state[194]),
        .w707(state[195]),
        .w708(state[196]),
        .w709(state[197]),
        .w710(state[198]),
        .w711(state[199]),
        .w712(state[200]),
        .w713(state[201]),
        .w714(state[202]),
        .w715(state[203]),
        .w716(state[204]),
        .w717(state[205]),
        .w718(state[206]),
        .w719(state[207]),
        .w720(state[208]),
        .w721(state[209]),
        .w722(state[210]),
        .w723(state[211]),
        .w724(state[212]),
        .w725(state[213]),
        .w726(state[214]),
        .w727(state[215]),
        .w728(state[216]),
        .w729(state[217]),
        .w730(state[218]),
        .w731(state[219]),
        .w732(state[220]),
        .w733(state[221]),
        .w734(state[222]),
        .w735(state[223]),
        .w736(state[224]),
        .w737(state[225]),
        .w738(state[226]),
        .w739(state[227]),
        .w740(state[228]),
        .w741(state[229]),
        .w742(state[230]),
        .w743(state[231]),
        .w744(state[232]),
        .w745(state[233]),
        .w746(state[234]),
        .w747(state[235]),
        .w748(state[236]),
        .w749(state[237]),
        .w750(state[238]),
        .w751(state[239]),
        .w752(state[240]),
        .w753(state[241]),
        .w754(state[242]),
        .w755(state[243]),
        .w756(state[244]),
        .w757(state[245]),
        .w758(state[246]),
        .w759(state[247]),
        .w760(state[248]),
        .w761(state[249]),
        .w762(state[250]),
        .w763(state[251]),
        .w764(state[252]),
        .w765(state[253]),
        .w766(state[254]),
        .w767(state[255]),
        .w135585(next_state[0]),
        .w135586(next_state[1]),
        .w135587(next_state[2]),
        .w135588(next_state[3]),
        .w135589(next_state[4]),
        .w135590(next_state[5]),
        .w135591(next_state[6]),
        .w135592(next_state[7]),
        .w135593(next_state[8]),
        .w135594(next_state[9]),
        .w135595(next_state[10]),
        .w135596(next_state[11]),
        .w135597(next_state[12]),
        .w135598(next_state[13]),
        .w135599(next_state[14]),
        .w135600(next_state[15]),
        .w135601(next_state[16]),
        .w135602(next_state[17]),
        .w135603(next_state[18]),
        .w135604(next_state[19]),
        .w135605(next_state[20]),
        .w135606(next_state[21]),
        .w135607(next_state[22]),
        .w135608(next_state[23]),
        .w135609(next_state[24]),
        .w135610(next_state[25]),
        .w135611(next_state[26]),
        .w135612(next_state[27]),
        .w135613(next_state[28]),
        .w135614(next_state[29]),
        .w135615(next_state[30]),
        .w135616(next_state[31]),
        .w135617(next_state[32]),
        .w135618(next_state[33]),
        .w135619(next_state[34]),
        .w135620(next_state[35]),
        .w135621(next_state[36]),
        .w135622(next_state[37]),
        .w135623(next_state[38]),
        .w135624(next_state[39]),
        .w135625(next_state[40]),
        .w135626(next_state[41]),
        .w135627(next_state[42]),
        .w135628(next_state[43]),
        .w135629(next_state[44]),
        .w135630(next_state[45]),
        .w135631(next_state[46]),
        .w135632(next_state[47]),
        .w135633(next_state[48]),
        .w135634(next_state[49]),
        .w135635(next_state[50]),
        .w135636(next_state[51]),
        .w135637(next_state[52]),
        .w135638(next_state[53]),
        .w135639(next_state[54]),
        .w135640(next_state[55]),
        .w135641(next_state[56]),
        .w135642(next_state[57]),
        .w135643(next_state[58]),
        .w135644(next_state[59]),
        .w135645(next_state[60]),
        .w135646(next_state[61]),
        .w135647(next_state[62]),
        .w135648(next_state[63]),
        .w135649(next_state[64]),
        .w135650(next_state[65]),
        .w135651(next_state[66]),
        .w135652(next_state[67]),
        .w135653(next_state[68]),
        .w135654(next_state[69]),
        .w135655(next_state[70]),
        .w135656(next_state[71]),
        .w135657(next_state[72]),
        .w135658(next_state[73]),
        .w135659(next_state[74]),
        .w135660(next_state[75]),
        .w135661(next_state[76]),
        .w135662(next_state[77]),
        .w135663(next_state[78]),
        .w135664(next_state[79]),
        .w135665(next_state[80]),
        .w135666(next_state[81]),
        .w135667(next_state[82]),
        .w135668(next_state[83]),
        .w135669(next_state[84]),
        .w135670(next_state[85]),
        .w135671(next_state[86]),
        .w135672(next_state[87]),
        .w135673(next_state[88]),
        .w135674(next_state[89]),
        .w135675(next_state[90]),
        .w135676(next_state[91]),
        .w135677(next_state[92]),
        .w135678(next_state[93]),
        .w135679(next_state[94]),
        .w135680(next_state[95]),
        .w135681(next_state[96]),
        .w135682(next_state[97]),
        .w135683(next_state[98]),
        .w135684(next_state[99]),
        .w135685(next_state[100]),
        .w135686(next_state[101]),
        .w135687(next_state[102]),
        .w135688(next_state[103]),
        .w135689(next_state[104]),
        .w135690(next_state[105]),
        .w135691(next_state[106]),
        .w135692(next_state[107]),
        .w135693(next_state[108]),
        .w135694(next_state[109]),
        .w135695(next_state[110]),
        .w135696(next_state[111]),
        .w135697(next_state[112]),
        .w135698(next_state[113]),
        .w135699(next_state[114]),
        .w135700(next_state[115]),
        .w135701(next_state[116]),
        .w135702(next_state[117]),
        .w135703(next_state[118]),
        .w135704(next_state[119]),
        .w135705(next_state[120]),
        .w135706(next_state[121]),
        .w135707(next_state[122]),
        .w135708(next_state[123]),
        .w135709(next_state[124]),
        .w135710(next_state[125]),
        .w135711(next_state[126]),
        .w135712(next_state[127]),
        .w135713(next_state[128]),
        .w135714(next_state[129]),
        .w135715(next_state[130]),
        .w135716(next_state[131]),
        .w135717(next_state[132]),
        .w135718(next_state[133]),
        .w135719(next_state[134]),
        .w135720(next_state[135]),
        .w135721(next_state[136]),
        .w135722(next_state[137]),
        .w135723(next_state[138]),
        .w135724(next_state[139]),
        .w135725(next_state[140]),
        .w135726(next_state[141]),
        .w135727(next_state[142]),
        .w135728(next_state[143]),
        .w135729(next_state[144]),
        .w135730(next_state[145]),
        .w135731(next_state[146]),
        .w135732(next_state[147]),
        .w135733(next_state[148]),
        .w135734(next_state[149]),
        .w135735(next_state[150]),
        .w135736(next_state[151]),
        .w135737(next_state[152]),
        .w135738(next_state[153]),
        .w135739(next_state[154]),
        .w135740(next_state[155]),
        .w135741(next_state[156]),
        .w135742(next_state[157]),
        .w135743(next_state[158]),
        .w135744(next_state[159]),
        .w135745(next_state[160]),
        .w135746(next_state[161]),
        .w135747(next_state[162]),
        .w135748(next_state[163]),
        .w135749(next_state[164]),
        .w135750(next_state[165]),
        .w135751(next_state[166]),
        .w135752(next_state[167]),
        .w135753(next_state[168]),
        .w135754(next_state[169]),
        .w135755(next_state[170]),
        .w135756(next_state[171]),
        .w135757(next_state[172]),
        .w135758(next_state[173]),
        .w135759(next_state[174]),
        .w135760(next_state[175]),
        .w135761(next_state[176]),
        .w135762(next_state[177]),
        .w135763(next_state[178]),
        .w135764(next_state[179]),
        .w135765(next_state[180]),
        .w135766(next_state[181]),
        .w135767(next_state[182]),
        .w135768(next_state[183]),
        .w135769(next_state[184]),
        .w135770(next_state[185]),
        .w135771(next_state[186]),
        .w135772(next_state[187]),
        .w135773(next_state[188]),
        .w135774(next_state[189]),
        .w135775(next_state[190]),
        .w135776(next_state[191]),
        .w135777(next_state[192]),
        .w135778(next_state[193]),
        .w135779(next_state[194]),
        .w135780(next_state[195]),
        .w135781(next_state[196]),
        .w135782(next_state[197]),
        .w135783(next_state[198]),
        .w135784(next_state[199]),
        .w135785(next_state[200]),
        .w135786(next_state[201]),
        .w135787(next_state[202]),
        .w135788(next_state[203]),
        .w135789(next_state[204]),
        .w135790(next_state[205]),
        .w135791(next_state[206]),
        .w135792(next_state[207]),
        .w135793(next_state[208]),
        .w135794(next_state[209]),
        .w135795(next_state[210]),
        .w135796(next_state[211]),
        .w135797(next_state[212]),
        .w135798(next_state[213]),
        .w135799(next_state[214]),
        .w135800(next_state[215]),
        .w135801(next_state[216]),
        .w135802(next_state[217]),
        .w135803(next_state[218]),
        .w135804(next_state[219]),
        .w135805(next_state[220]),
        .w135806(next_state[221]),
        .w135807(next_state[222]),
        .w135808(next_state[223]),
        .w135809(next_state[224]),
        .w135810(next_state[225]),
        .w135811(next_state[226]),
        .w135812(next_state[227]),
        .w135813(next_state[228]),
        .w135814(next_state[229]),
        .w135815(next_state[230]),
        .w135816(next_state[231]),
        .w135817(next_state[232]),
        .w135818(next_state[233]),
        .w135819(next_state[234]),
        .w135820(next_state[235]),
        .w135821(next_state[236]),
        .w135822(next_state[237]),
        .w135823(next_state[238]),
        .w135824(next_state[239]),
        .w135825(next_state[240]),
        .w135826(next_state[241]),
        .w135827(next_state[242]),
        .w135828(next_state[243]),
        .w135829(next_state[244]),
        .w135830(next_state[245]),
        .w135831(next_state[246]),
        .w135832(next_state[247]),
        .w135833(next_state[248]),
        .w135834(next_state[249]),
        .w135835(next_state[250]),
        .w135836(next_state[251]),
        .w135837(next_state[252]),
        .w135838(next_state[253]),
        .w135839(next_state[254]),
        .w135840(next_state[255]),
);
endmodule